
`timescale 1ns / 1ps
module cache_tb();

localparam INDEX_WIDTH          = 3;
localparam WORD_OFFSET_WIDTH    = 1;
localparam TOTAL_WORD_NUM       = 1024;

// cache test
reg [31:0]  i_addr_rom [TOTAL_WORD_NUM];
reg [31:0]  d_addr_rom [TOTAL_WORD_NUM];
reg [31:0]  data_ram [TOTAL_WORD_NUM];
reg         wvalid_rom [TOTAL_WORD_NUM];
reg [31:0]  wdata_rom [TOTAL_WORD_NUM];
reg [31:0]  i_test_index = 0;
reg [31:0]  d_test_index = 0;
reg clk = 1'b1, rstn = 1'b0;

initial #5 rstn = 1'b1; 
always #1 clk = ~clk;

// generate data_ram
initial begin
    data_ram[    0] = 'h00000000; 	    data_ram[    1] = 'h00000001; 	    data_ram[    2] = 'h00000002; 	    data_ram[    3] = 'h00000003; 	    data_ram[    4] = 'h00000004; 	    data_ram[    5] = 'h00000005; 	    data_ram[    6] = 'h00000006; 	    data_ram[    7] = 'h00000007; 	
    data_ram[    8] = 'h00000008; 	    data_ram[    9] = 'h00000009; 	    data_ram[   10] = 'h0000000a; 	    data_ram[   11] = 'h0000000b; 	    data_ram[   12] = 'h0000000c; 	    data_ram[   13] = 'h0000000d; 	    data_ram[   14] = 'h0000000e; 	    data_ram[   15] = 'h0000000f; 	
    data_ram[   16] = 'h00000010; 	    data_ram[   17] = 'h00000011; 	    data_ram[   18] = 'h00000012; 	    data_ram[   19] = 'h00000013; 	    data_ram[   20] = 'h00000014; 	    data_ram[   21] = 'h00000015; 	    data_ram[   22] = 'h00000016; 	    data_ram[   23] = 'h00000017; 	
    data_ram[   24] = 'h00000018; 	    data_ram[   25] = 'h00000019; 	    data_ram[   26] = 'h0000001a; 	    data_ram[   27] = 'h0000001b; 	    data_ram[   28] = 'h0000001c; 	    data_ram[   29] = 'h0000001d; 	    data_ram[   30] = 'h0000001e; 	    data_ram[   31] = 'h0000001f; 	
    data_ram[   32] = 'h00000020; 	    data_ram[   33] = 'h00000021; 	    data_ram[   34] = 'h00000022; 	    data_ram[   35] = 'h00000023; 	    data_ram[   36] = 'h00000024; 	    data_ram[   37] = 'h00000025; 	    data_ram[   38] = 'h00000026; 	    data_ram[   39] = 'h00000027; 	
    data_ram[   40] = 'h00000028; 	    data_ram[   41] = 'h00000029; 	    data_ram[   42] = 'h0000002a; 	    data_ram[   43] = 'h0000002b; 	    data_ram[   44] = 'h0000002c; 	    data_ram[   45] = 'h0000002d; 	    data_ram[   46] = 'h0000002e; 	    data_ram[   47] = 'h0000002f; 	
    data_ram[   48] = 'h00000030; 	    data_ram[   49] = 'h00000031; 	    data_ram[   50] = 'h00000032; 	    data_ram[   51] = 'h00000033; 	    data_ram[   52] = 'h00000034; 	    data_ram[   53] = 'h00000035; 	    data_ram[   54] = 'h00000036; 	    data_ram[   55] = 'h00000037; 	
    data_ram[   56] = 'h00000038; 	    data_ram[   57] = 'h00000039; 	    data_ram[   58] = 'h0000003a; 	    data_ram[   59] = 'h0000003b; 	    data_ram[   60] = 'h0000003c; 	    data_ram[   61] = 'h0000003d; 	    data_ram[   62] = 'h0000003e; 	    data_ram[   63] = 'h0000003f; 	
    data_ram[   64] = 'h00000040; 	    data_ram[   65] = 'h00000041; 	    data_ram[   66] = 'h00000042; 	    data_ram[   67] = 'h00000043; 	    data_ram[   68] = 'h00000044; 	    data_ram[   69] = 'h00000045; 	    data_ram[   70] = 'h00000046; 	    data_ram[   71] = 'h00000047; 	
    data_ram[   72] = 'h00000048; 	    data_ram[   73] = 'h00000049; 	    data_ram[   74] = 'h0000004a; 	    data_ram[   75] = 'h0000004b; 	    data_ram[   76] = 'h0000004c; 	    data_ram[   77] = 'h0000004d; 	    data_ram[   78] = 'h0000004e; 	    data_ram[   79] = 'h0000004f; 	
    data_ram[   80] = 'h00000050; 	    data_ram[   81] = 'h00000051; 	    data_ram[   82] = 'h00000052; 	    data_ram[   83] = 'h00000053; 	    data_ram[   84] = 'h00000054; 	    data_ram[   85] = 'h00000055; 	    data_ram[   86] = 'h00000056; 	    data_ram[   87] = 'h00000057; 	
    data_ram[   88] = 'h00000058; 	    data_ram[   89] = 'h00000059; 	    data_ram[   90] = 'h0000005a; 	    data_ram[   91] = 'h0000005b; 	    data_ram[   92] = 'h0000005c; 	    data_ram[   93] = 'h0000005d; 	    data_ram[   94] = 'h0000005e; 	    data_ram[   95] = 'h0000005f; 	
    data_ram[   96] = 'h00000060; 	    data_ram[   97] = 'h00000061; 	    data_ram[   98] = 'h00000062; 	    data_ram[   99] = 'h00000063; 	    data_ram[  100] = 'h00000064; 	    data_ram[  101] = 'h00000065; 	    data_ram[  102] = 'h00000066; 	    data_ram[  103] = 'h00000067; 	
    data_ram[  104] = 'h00000068; 	    data_ram[  105] = 'h00000069; 	    data_ram[  106] = 'h0000006a; 	    data_ram[  107] = 'h0000006b; 	    data_ram[  108] = 'h0000006c; 	    data_ram[  109] = 'h0000006d; 	    data_ram[  110] = 'h0000006e; 	    data_ram[  111] = 'h0000006f; 	
    data_ram[  112] = 'h00000070; 	    data_ram[  113] = 'h00000071; 	    data_ram[  114] = 'h00000072; 	    data_ram[  115] = 'h00000073; 	    data_ram[  116] = 'h00000074; 	    data_ram[  117] = 'h00000075; 	    data_ram[  118] = 'h00000076; 	    data_ram[  119] = 'h00000077; 	
    data_ram[  120] = 'h00000078; 	    data_ram[  121] = 'h00000079; 	    data_ram[  122] = 'h0000007a; 	    data_ram[  123] = 'h0000007b; 	    data_ram[  124] = 'h0000007c; 	    data_ram[  125] = 'h0000007d; 	    data_ram[  126] = 'h0000007e; 	    data_ram[  127] = 'h0000007f; 	
    data_ram[  128] = 'h00000080; 	    data_ram[  129] = 'h00000081; 	    data_ram[  130] = 'h00000082; 	    data_ram[  131] = 'h00000083; 	    data_ram[  132] = 'h00000084; 	    data_ram[  133] = 'h00000085; 	    data_ram[  134] = 'h00000086; 	    data_ram[  135] = 'h00000087; 	
    data_ram[  136] = 'h00000088; 	    data_ram[  137] = 'h00000089; 	    data_ram[  138] = 'h0000008a; 	    data_ram[  139] = 'h0000008b; 	    data_ram[  140] = 'h0000008c; 	    data_ram[  141] = 'h0000008d; 	    data_ram[  142] = 'h0000008e; 	    data_ram[  143] = 'h0000008f; 	
    data_ram[  144] = 'h00000090; 	    data_ram[  145] = 'h00000091; 	    data_ram[  146] = 'h00000092; 	    data_ram[  147] = 'h00000093; 	    data_ram[  148] = 'h00000094; 	    data_ram[  149] = 'h00000095; 	    data_ram[  150] = 'h00000096; 	    data_ram[  151] = 'h00000097; 	
    data_ram[  152] = 'h00000098; 	    data_ram[  153] = 'h00000099; 	    data_ram[  154] = 'h0000009a; 	    data_ram[  155] = 'h0000009b; 	    data_ram[  156] = 'h0000009c; 	    data_ram[  157] = 'h0000009d; 	    data_ram[  158] = 'h0000009e; 	    data_ram[  159] = 'h0000009f; 	
    data_ram[  160] = 'h000000a0; 	    data_ram[  161] = 'h000000a1; 	    data_ram[  162] = 'h000000a2; 	    data_ram[  163] = 'h000000a3; 	    data_ram[  164] = 'h000000a4; 	    data_ram[  165] = 'h000000a5; 	    data_ram[  166] = 'h000000a6; 	    data_ram[  167] = 'h000000a7; 	
    data_ram[  168] = 'h000000a8; 	    data_ram[  169] = 'h000000a9; 	    data_ram[  170] = 'h000000aa; 	    data_ram[  171] = 'h000000ab; 	    data_ram[  172] = 'h000000ac; 	    data_ram[  173] = 'h000000ad; 	    data_ram[  174] = 'h000000ae; 	    data_ram[  175] = 'h000000af; 	
    data_ram[  176] = 'h000000b0; 	    data_ram[  177] = 'h000000b1; 	    data_ram[  178] = 'h000000b2; 	    data_ram[  179] = 'h000000b3; 	    data_ram[  180] = 'h000000b4; 	    data_ram[  181] = 'h000000b5; 	    data_ram[  182] = 'h000000b6; 	    data_ram[  183] = 'h000000b7; 	
    data_ram[  184] = 'h000000b8; 	    data_ram[  185] = 'h000000b9; 	    data_ram[  186] = 'h000000ba; 	    data_ram[  187] = 'h000000bb; 	    data_ram[  188] = 'h000000bc; 	    data_ram[  189] = 'h000000bd; 	    data_ram[  190] = 'h000000be; 	    data_ram[  191] = 'h000000bf; 	
    data_ram[  192] = 'h000000c0; 	    data_ram[  193] = 'h000000c1; 	    data_ram[  194] = 'h000000c2; 	    data_ram[  195] = 'h000000c3; 	    data_ram[  196] = 'h000000c4; 	    data_ram[  197] = 'h000000c5; 	    data_ram[  198] = 'h000000c6; 	    data_ram[  199] = 'h000000c7; 	
    data_ram[  200] = 'h000000c8; 	    data_ram[  201] = 'h000000c9; 	    data_ram[  202] = 'h000000ca; 	    data_ram[  203] = 'h000000cb; 	    data_ram[  204] = 'h000000cc; 	    data_ram[  205] = 'h000000cd; 	    data_ram[  206] = 'h000000ce; 	    data_ram[  207] = 'h000000cf; 	
    data_ram[  208] = 'h000000d0; 	    data_ram[  209] = 'h000000d1; 	    data_ram[  210] = 'h000000d2; 	    data_ram[  211] = 'h000000d3; 	    data_ram[  212] = 'h000000d4; 	    data_ram[  213] = 'h000000d5; 	    data_ram[  214] = 'h000000d6; 	    data_ram[  215] = 'h000000d7; 	
    data_ram[  216] = 'h000000d8; 	    data_ram[  217] = 'h000000d9; 	    data_ram[  218] = 'h000000da; 	    data_ram[  219] = 'h000000db; 	    data_ram[  220] = 'h000000dc; 	    data_ram[  221] = 'h000000dd; 	    data_ram[  222] = 'h000000de; 	    data_ram[  223] = 'h000000df; 	
    data_ram[  224] = 'h000000e0; 	    data_ram[  225] = 'h000000e1; 	    data_ram[  226] = 'h000000e2; 	    data_ram[  227] = 'h000000e3; 	    data_ram[  228] = 'h000000e4; 	    data_ram[  229] = 'h000000e5; 	    data_ram[  230] = 'h000000e6; 	    data_ram[  231] = 'h000000e7; 	
    data_ram[  232] = 'h000000e8; 	    data_ram[  233] = 'h000000e9; 	    data_ram[  234] = 'h000000ea; 	    data_ram[  235] = 'h000000eb; 	    data_ram[  236] = 'h000000ec; 	    data_ram[  237] = 'h000000ed; 	    data_ram[  238] = 'h000000ee; 	    data_ram[  239] = 'h000000ef; 	
    data_ram[  240] = 'h000000f0; 	    data_ram[  241] = 'h000000f1; 	    data_ram[  242] = 'h000000f2; 	    data_ram[  243] = 'h000000f3; 	    data_ram[  244] = 'h000000f4; 	    data_ram[  245] = 'h000000f5; 	    data_ram[  246] = 'h000000f6; 	    data_ram[  247] = 'h000000f7; 	
    data_ram[  248] = 'h000000f8; 	    data_ram[  249] = 'h000000f9; 	    data_ram[  250] = 'h000000fa; 	    data_ram[  251] = 'h000000fb; 	    data_ram[  252] = 'h000000fc; 	    data_ram[  253] = 'h000000fd; 	    data_ram[  254] = 'h000000fe; 	    data_ram[  255] = 'h000000ff; 	
    data_ram[  256] = 'h00000100; 	    data_ram[  257] = 'h00000101; 	    data_ram[  258] = 'h00000102; 	    data_ram[  259] = 'h00000103; 	    data_ram[  260] = 'h00000104; 	    data_ram[  261] = 'h00000105; 	    data_ram[  262] = 'h00000106; 	    data_ram[  263] = 'h00000107; 	
    data_ram[  264] = 'h00000108; 	    data_ram[  265] = 'h00000109; 	    data_ram[  266] = 'h0000010a; 	    data_ram[  267] = 'h0000010b; 	    data_ram[  268] = 'h0000010c; 	    data_ram[  269] = 'h0000010d; 	    data_ram[  270] = 'h0000010e; 	    data_ram[  271] = 'h0000010f; 	
    data_ram[  272] = 'h00000110; 	    data_ram[  273] = 'h00000111; 	    data_ram[  274] = 'h00000112; 	    data_ram[  275] = 'h00000113; 	    data_ram[  276] = 'h00000114; 	    data_ram[  277] = 'h00000115; 	    data_ram[  278] = 'h00000116; 	    data_ram[  279] = 'h00000117; 	
    data_ram[  280] = 'h00000118; 	    data_ram[  281] = 'h00000119; 	    data_ram[  282] = 'h0000011a; 	    data_ram[  283] = 'h0000011b; 	    data_ram[  284] = 'h0000011c; 	    data_ram[  285] = 'h0000011d; 	    data_ram[  286] = 'h0000011e; 	    data_ram[  287] = 'h0000011f; 	
    data_ram[  288] = 'h00000120; 	    data_ram[  289] = 'h00000121; 	    data_ram[  290] = 'h00000122; 	    data_ram[  291] = 'h00000123; 	    data_ram[  292] = 'h00000124; 	    data_ram[  293] = 'h00000125; 	    data_ram[  294] = 'h00000126; 	    data_ram[  295] = 'h00000127; 	
    data_ram[  296] = 'h00000128; 	    data_ram[  297] = 'h00000129; 	    data_ram[  298] = 'h0000012a; 	    data_ram[  299] = 'h0000012b; 	    data_ram[  300] = 'h0000012c; 	    data_ram[  301] = 'h0000012d; 	    data_ram[  302] = 'h0000012e; 	    data_ram[  303] = 'h0000012f; 	
    data_ram[  304] = 'h00000130; 	    data_ram[  305] = 'h00000131; 	    data_ram[  306] = 'h00000132; 	    data_ram[  307] = 'h00000133; 	    data_ram[  308] = 'h00000134; 	    data_ram[  309] = 'h00000135; 	    data_ram[  310] = 'h00000136; 	    data_ram[  311] = 'h00000137; 	
    data_ram[  312] = 'h00000138; 	    data_ram[  313] = 'h00000139; 	    data_ram[  314] = 'h0000013a; 	    data_ram[  315] = 'h0000013b; 	    data_ram[  316] = 'h0000013c; 	    data_ram[  317] = 'h0000013d; 	    data_ram[  318] = 'h0000013e; 	    data_ram[  319] = 'h0000013f; 	
    data_ram[  320] = 'h00000140; 	    data_ram[  321] = 'h00000141; 	    data_ram[  322] = 'h00000142; 	    data_ram[  323] = 'h00000143; 	    data_ram[  324] = 'h00000144; 	    data_ram[  325] = 'h00000145; 	    data_ram[  326] = 'h00000146; 	    data_ram[  327] = 'h00000147; 	
    data_ram[  328] = 'h00000148; 	    data_ram[  329] = 'h00000149; 	    data_ram[  330] = 'h0000014a; 	    data_ram[  331] = 'h0000014b; 	    data_ram[  332] = 'h0000014c; 	    data_ram[  333] = 'h0000014d; 	    data_ram[  334] = 'h0000014e; 	    data_ram[  335] = 'h0000014f; 	
    data_ram[  336] = 'h00000150; 	    data_ram[  337] = 'h00000151; 	    data_ram[  338] = 'h00000152; 	    data_ram[  339] = 'h00000153; 	    data_ram[  340] = 'h00000154; 	    data_ram[  341] = 'h00000155; 	    data_ram[  342] = 'h00000156; 	    data_ram[  343] = 'h00000157; 	
    data_ram[  344] = 'h00000158; 	    data_ram[  345] = 'h00000159; 	    data_ram[  346] = 'h0000015a; 	    data_ram[  347] = 'h0000015b; 	    data_ram[  348] = 'h0000015c; 	    data_ram[  349] = 'h0000015d; 	    data_ram[  350] = 'h0000015e; 	    data_ram[  351] = 'h0000015f; 	
    data_ram[  352] = 'h00000160; 	    data_ram[  353] = 'h00000161; 	    data_ram[  354] = 'h00000162; 	    data_ram[  355] = 'h00000163; 	    data_ram[  356] = 'h00000164; 	    data_ram[  357] = 'h00000165; 	    data_ram[  358] = 'h00000166; 	    data_ram[  359] = 'h00000167; 	
    data_ram[  360] = 'h00000168; 	    data_ram[  361] = 'h00000169; 	    data_ram[  362] = 'h0000016a; 	    data_ram[  363] = 'h0000016b; 	    data_ram[  364] = 'h0000016c; 	    data_ram[  365] = 'h0000016d; 	    data_ram[  366] = 'h0000016e; 	    data_ram[  367] = 'h0000016f; 	
    data_ram[  368] = 'h00000170; 	    data_ram[  369] = 'h00000171; 	    data_ram[  370] = 'h00000172; 	    data_ram[  371] = 'h00000173; 	    data_ram[  372] = 'h00000174; 	    data_ram[  373] = 'h00000175; 	    data_ram[  374] = 'h00000176; 	    data_ram[  375] = 'h00000177; 	
    data_ram[  376] = 'h00000178; 	    data_ram[  377] = 'h00000179; 	    data_ram[  378] = 'h0000017a; 	    data_ram[  379] = 'h0000017b; 	    data_ram[  380] = 'h0000017c; 	    data_ram[  381] = 'h0000017d; 	    data_ram[  382] = 'h0000017e; 	    data_ram[  383] = 'h0000017f; 	
    data_ram[  384] = 'h00000180; 	    data_ram[  385] = 'h00000181; 	    data_ram[  386] = 'h00000182; 	    data_ram[  387] = 'h00000183; 	    data_ram[  388] = 'h00000184; 	    data_ram[  389] = 'h00000185; 	    data_ram[  390] = 'h00000186; 	    data_ram[  391] = 'h00000187; 	
    data_ram[  392] = 'h00000188; 	    data_ram[  393] = 'h00000189; 	    data_ram[  394] = 'h0000018a; 	    data_ram[  395] = 'h0000018b; 	    data_ram[  396] = 'h0000018c; 	    data_ram[  397] = 'h0000018d; 	    data_ram[  398] = 'h0000018e; 	    data_ram[  399] = 'h0000018f; 	
    data_ram[  400] = 'h00000190; 	    data_ram[  401] = 'h00000191; 	    data_ram[  402] = 'h00000192; 	    data_ram[  403] = 'h00000193; 	    data_ram[  404] = 'h00000194; 	    data_ram[  405] = 'h00000195; 	    data_ram[  406] = 'h00000196; 	    data_ram[  407] = 'h00000197; 	
    data_ram[  408] = 'h00000198; 	    data_ram[  409] = 'h00000199; 	    data_ram[  410] = 'h0000019a; 	    data_ram[  411] = 'h0000019b; 	    data_ram[  412] = 'h0000019c; 	    data_ram[  413] = 'h0000019d; 	    data_ram[  414] = 'h0000019e; 	    data_ram[  415] = 'h0000019f; 	
    data_ram[  416] = 'h000001a0; 	    data_ram[  417] = 'h000001a1; 	    data_ram[  418] = 'h000001a2; 	    data_ram[  419] = 'h000001a3; 	    data_ram[  420] = 'h000001a4; 	    data_ram[  421] = 'h000001a5; 	    data_ram[  422] = 'h000001a6; 	    data_ram[  423] = 'h000001a7; 	
    data_ram[  424] = 'h000001a8; 	    data_ram[  425] = 'h000001a9; 	    data_ram[  426] = 'h000001aa; 	    data_ram[  427] = 'h000001ab; 	    data_ram[  428] = 'h000001ac; 	    data_ram[  429] = 'h000001ad; 	    data_ram[  430] = 'h000001ae; 	    data_ram[  431] = 'h000001af; 	
    data_ram[  432] = 'h000001b0; 	    data_ram[  433] = 'h000001b1; 	    data_ram[  434] = 'h000001b2; 	    data_ram[  435] = 'h000001b3; 	    data_ram[  436] = 'h000001b4; 	    data_ram[  437] = 'h000001b5; 	    data_ram[  438] = 'h000001b6; 	    data_ram[  439] = 'h000001b7; 	
    data_ram[  440] = 'h000001b8; 	    data_ram[  441] = 'h000001b9; 	    data_ram[  442] = 'h000001ba; 	    data_ram[  443] = 'h000001bb; 	    data_ram[  444] = 'h000001bc; 	    data_ram[  445] = 'h000001bd; 	    data_ram[  446] = 'h000001be; 	    data_ram[  447] = 'h000001bf; 	
    data_ram[  448] = 'h000001c0; 	    data_ram[  449] = 'h000001c1; 	    data_ram[  450] = 'h000001c2; 	    data_ram[  451] = 'h000001c3; 	    data_ram[  452] = 'h000001c4; 	    data_ram[  453] = 'h000001c5; 	    data_ram[  454] = 'h000001c6; 	    data_ram[  455] = 'h000001c7; 	
    data_ram[  456] = 'h000001c8; 	    data_ram[  457] = 'h000001c9; 	    data_ram[  458] = 'h000001ca; 	    data_ram[  459] = 'h000001cb; 	    data_ram[  460] = 'h000001cc; 	    data_ram[  461] = 'h000001cd; 	    data_ram[  462] = 'h000001ce; 	    data_ram[  463] = 'h000001cf; 	
    data_ram[  464] = 'h000001d0; 	    data_ram[  465] = 'h000001d1; 	    data_ram[  466] = 'h000001d2; 	    data_ram[  467] = 'h000001d3; 	    data_ram[  468] = 'h000001d4; 	    data_ram[  469] = 'h000001d5; 	    data_ram[  470] = 'h000001d6; 	    data_ram[  471] = 'h000001d7; 	
    data_ram[  472] = 'h000001d8; 	    data_ram[  473] = 'h000001d9; 	    data_ram[  474] = 'h000001da; 	    data_ram[  475] = 'h000001db; 	    data_ram[  476] = 'h000001dc; 	    data_ram[  477] = 'h000001dd; 	    data_ram[  478] = 'h000001de; 	    data_ram[  479] = 'h000001df; 	
    data_ram[  480] = 'h000001e0; 	    data_ram[  481] = 'h000001e1; 	    data_ram[  482] = 'h000001e2; 	    data_ram[  483] = 'h000001e3; 	    data_ram[  484] = 'h000001e4; 	    data_ram[  485] = 'h000001e5; 	    data_ram[  486] = 'h000001e6; 	    data_ram[  487] = 'h000001e7; 	
    data_ram[  488] = 'h000001e8; 	    data_ram[  489] = 'h000001e9; 	    data_ram[  490] = 'h000001ea; 	    data_ram[  491] = 'h000001eb; 	    data_ram[  492] = 'h000001ec; 	    data_ram[  493] = 'h000001ed; 	    data_ram[  494] = 'h000001ee; 	    data_ram[  495] = 'h000001ef; 	
    data_ram[  496] = 'h000001f0; 	    data_ram[  497] = 'h000001f1; 	    data_ram[  498] = 'h000001f2; 	    data_ram[  499] = 'h000001f3; 	    data_ram[  500] = 'h000001f4; 	    data_ram[  501] = 'h000001f5; 	    data_ram[  502] = 'h000001f6; 	    data_ram[  503] = 'h000001f7; 	
    data_ram[  504] = 'h000001f8; 	    data_ram[  505] = 'h000001f9; 	    data_ram[  506] = 'h000001fa; 	    data_ram[  507] = 'h000001fb; 	    data_ram[  508] = 'h000001fc; 	    data_ram[  509] = 'h000001fd; 	    data_ram[  510] = 'h000001fe; 	    data_ram[  511] = 'h000001ff; 	
    data_ram[  512] = 'h00000200; 	    data_ram[  513] = 'h00000201; 	    data_ram[  514] = 'h00000202; 	    data_ram[  515] = 'h00000203; 	    data_ram[  516] = 'h00000204; 	    data_ram[  517] = 'h00000205; 	    data_ram[  518] = 'h00000206; 	    data_ram[  519] = 'h00000207; 	
    data_ram[  520] = 'h00000208; 	    data_ram[  521] = 'h00000209; 	    data_ram[  522] = 'h0000020a; 	    data_ram[  523] = 'h0000020b; 	    data_ram[  524] = 'h0000020c; 	    data_ram[  525] = 'h0000020d; 	    data_ram[  526] = 'h0000020e; 	    data_ram[  527] = 'h0000020f; 	
    data_ram[  528] = 'h00000210; 	    data_ram[  529] = 'h00000211; 	    data_ram[  530] = 'h00000212; 	    data_ram[  531] = 'h00000213; 	    data_ram[  532] = 'h00000214; 	    data_ram[  533] = 'h00000215; 	    data_ram[  534] = 'h00000216; 	    data_ram[  535] = 'h00000217; 	
    data_ram[  536] = 'h00000218; 	    data_ram[  537] = 'h00000219; 	    data_ram[  538] = 'h0000021a; 	    data_ram[  539] = 'h0000021b; 	    data_ram[  540] = 'h0000021c; 	    data_ram[  541] = 'h0000021d; 	    data_ram[  542] = 'h0000021e; 	    data_ram[  543] = 'h0000021f; 	
    data_ram[  544] = 'h00000220; 	    data_ram[  545] = 'h00000221; 	    data_ram[  546] = 'h00000222; 	    data_ram[  547] = 'h00000223; 	    data_ram[  548] = 'h00000224; 	    data_ram[  549] = 'h00000225; 	    data_ram[  550] = 'h00000226; 	    data_ram[  551] = 'h00000227; 	
    data_ram[  552] = 'h00000228; 	    data_ram[  553] = 'h00000229; 	    data_ram[  554] = 'h0000022a; 	    data_ram[  555] = 'h0000022b; 	    data_ram[  556] = 'h0000022c; 	    data_ram[  557] = 'h0000022d; 	    data_ram[  558] = 'h0000022e; 	    data_ram[  559] = 'h0000022f; 	
    data_ram[  560] = 'h00000230; 	    data_ram[  561] = 'h00000231; 	    data_ram[  562] = 'h00000232; 	    data_ram[  563] = 'h00000233; 	    data_ram[  564] = 'h00000234; 	    data_ram[  565] = 'h00000235; 	    data_ram[  566] = 'h00000236; 	    data_ram[  567] = 'h00000237; 	
    data_ram[  568] = 'h00000238; 	    data_ram[  569] = 'h00000239; 	    data_ram[  570] = 'h0000023a; 	    data_ram[  571] = 'h0000023b; 	    data_ram[  572] = 'h0000023c; 	    data_ram[  573] = 'h0000023d; 	    data_ram[  574] = 'h0000023e; 	    data_ram[  575] = 'h0000023f; 	
    data_ram[  576] = 'h00000240; 	    data_ram[  577] = 'h00000241; 	    data_ram[  578] = 'h00000242; 	    data_ram[  579] = 'h00000243; 	    data_ram[  580] = 'h00000244; 	    data_ram[  581] = 'h00000245; 	    data_ram[  582] = 'h00000246; 	    data_ram[  583] = 'h00000247; 	
    data_ram[  584] = 'h00000248; 	    data_ram[  585] = 'h00000249; 	    data_ram[  586] = 'h0000024a; 	    data_ram[  587] = 'h0000024b; 	    data_ram[  588] = 'h0000024c; 	    data_ram[  589] = 'h0000024d; 	    data_ram[  590] = 'h0000024e; 	    data_ram[  591] = 'h0000024f; 	
    data_ram[  592] = 'h00000250; 	    data_ram[  593] = 'h00000251; 	    data_ram[  594] = 'h00000252; 	    data_ram[  595] = 'h00000253; 	    data_ram[  596] = 'h00000254; 	    data_ram[  597] = 'h00000255; 	    data_ram[  598] = 'h00000256; 	    data_ram[  599] = 'h00000257; 	
    data_ram[  600] = 'h00000258; 	    data_ram[  601] = 'h00000259; 	    data_ram[  602] = 'h0000025a; 	    data_ram[  603] = 'h0000025b; 	    data_ram[  604] = 'h0000025c; 	    data_ram[  605] = 'h0000025d; 	    data_ram[  606] = 'h0000025e; 	    data_ram[  607] = 'h0000025f; 	
    data_ram[  608] = 'h00000260; 	    data_ram[  609] = 'h00000261; 	    data_ram[  610] = 'h00000262; 	    data_ram[  611] = 'h00000263; 	    data_ram[  612] = 'h00000264; 	    data_ram[  613] = 'h00000265; 	    data_ram[  614] = 'h00000266; 	    data_ram[  615] = 'h00000267; 	
    data_ram[  616] = 'h00000268; 	    data_ram[  617] = 'h00000269; 	    data_ram[  618] = 'h0000026a; 	    data_ram[  619] = 'h0000026b; 	    data_ram[  620] = 'h0000026c; 	    data_ram[  621] = 'h0000026d; 	    data_ram[  622] = 'h0000026e; 	    data_ram[  623] = 'h0000026f; 	
    data_ram[  624] = 'h00000270; 	    data_ram[  625] = 'h00000271; 	    data_ram[  626] = 'h00000272; 	    data_ram[  627] = 'h00000273; 	    data_ram[  628] = 'h00000274; 	    data_ram[  629] = 'h00000275; 	    data_ram[  630] = 'h00000276; 	    data_ram[  631] = 'h00000277; 	
    data_ram[  632] = 'h00000278; 	    data_ram[  633] = 'h00000279; 	    data_ram[  634] = 'h0000027a; 	    data_ram[  635] = 'h0000027b; 	    data_ram[  636] = 'h0000027c; 	    data_ram[  637] = 'h0000027d; 	    data_ram[  638] = 'h0000027e; 	    data_ram[  639] = 'h0000027f; 	
    data_ram[  640] = 'h00000280; 	    data_ram[  641] = 'h00000281; 	    data_ram[  642] = 'h00000282; 	    data_ram[  643] = 'h00000283; 	    data_ram[  644] = 'h00000284; 	    data_ram[  645] = 'h00000285; 	    data_ram[  646] = 'h00000286; 	    data_ram[  647] = 'h00000287; 	
    data_ram[  648] = 'h00000288; 	    data_ram[  649] = 'h00000289; 	    data_ram[  650] = 'h0000028a; 	    data_ram[  651] = 'h0000028b; 	    data_ram[  652] = 'h0000028c; 	    data_ram[  653] = 'h0000028d; 	    data_ram[  654] = 'h0000028e; 	    data_ram[  655] = 'h0000028f; 	
    data_ram[  656] = 'h00000290; 	    data_ram[  657] = 'h00000291; 	    data_ram[  658] = 'h00000292; 	    data_ram[  659] = 'h00000293; 	    data_ram[  660] = 'h00000294; 	    data_ram[  661] = 'h00000295; 	    data_ram[  662] = 'h00000296; 	    data_ram[  663] = 'h00000297; 	
    data_ram[  664] = 'h00000298; 	    data_ram[  665] = 'h00000299; 	    data_ram[  666] = 'h0000029a; 	    data_ram[  667] = 'h0000029b; 	    data_ram[  668] = 'h0000029c; 	    data_ram[  669] = 'h0000029d; 	    data_ram[  670] = 'h0000029e; 	    data_ram[  671] = 'h0000029f; 	
    data_ram[  672] = 'h000002a0; 	    data_ram[  673] = 'h000002a1; 	    data_ram[  674] = 'h000002a2; 	    data_ram[  675] = 'h000002a3; 	    data_ram[  676] = 'h000002a4; 	    data_ram[  677] = 'h000002a5; 	    data_ram[  678] = 'h000002a6; 	    data_ram[  679] = 'h000002a7; 	
    data_ram[  680] = 'h000002a8; 	    data_ram[  681] = 'h000002a9; 	    data_ram[  682] = 'h000002aa; 	    data_ram[  683] = 'h000002ab; 	    data_ram[  684] = 'h000002ac; 	    data_ram[  685] = 'h000002ad; 	    data_ram[  686] = 'h000002ae; 	    data_ram[  687] = 'h000002af; 	
    data_ram[  688] = 'h000002b0; 	    data_ram[  689] = 'h000002b1; 	    data_ram[  690] = 'h000002b2; 	    data_ram[  691] = 'h000002b3; 	    data_ram[  692] = 'h000002b4; 	    data_ram[  693] = 'h000002b5; 	    data_ram[  694] = 'h000002b6; 	    data_ram[  695] = 'h000002b7; 	
    data_ram[  696] = 'h000002b8; 	    data_ram[  697] = 'h000002b9; 	    data_ram[  698] = 'h000002ba; 	    data_ram[  699] = 'h000002bb; 	    data_ram[  700] = 'h000002bc; 	    data_ram[  701] = 'h000002bd; 	    data_ram[  702] = 'h000002be; 	    data_ram[  703] = 'h000002bf; 	
    data_ram[  704] = 'h000002c0; 	    data_ram[  705] = 'h000002c1; 	    data_ram[  706] = 'h000002c2; 	    data_ram[  707] = 'h000002c3; 	    data_ram[  708] = 'h000002c4; 	    data_ram[  709] = 'h000002c5; 	    data_ram[  710] = 'h000002c6; 	    data_ram[  711] = 'h000002c7; 	
    data_ram[  712] = 'h000002c8; 	    data_ram[  713] = 'h000002c9; 	    data_ram[  714] = 'h000002ca; 	    data_ram[  715] = 'h000002cb; 	    data_ram[  716] = 'h000002cc; 	    data_ram[  717] = 'h000002cd; 	    data_ram[  718] = 'h000002ce; 	    data_ram[  719] = 'h000002cf; 	
    data_ram[  720] = 'h000002d0; 	    data_ram[  721] = 'h000002d1; 	    data_ram[  722] = 'h000002d2; 	    data_ram[  723] = 'h000002d3; 	    data_ram[  724] = 'h000002d4; 	    data_ram[  725] = 'h000002d5; 	    data_ram[  726] = 'h000002d6; 	    data_ram[  727] = 'h000002d7; 	
    data_ram[  728] = 'h000002d8; 	    data_ram[  729] = 'h000002d9; 	    data_ram[  730] = 'h000002da; 	    data_ram[  731] = 'h000002db; 	    data_ram[  732] = 'h000002dc; 	    data_ram[  733] = 'h000002dd; 	    data_ram[  734] = 'h000002de; 	    data_ram[  735] = 'h000002df; 	
    data_ram[  736] = 'h000002e0; 	    data_ram[  737] = 'h000002e1; 	    data_ram[  738] = 'h000002e2; 	    data_ram[  739] = 'h000002e3; 	    data_ram[  740] = 'h000002e4; 	    data_ram[  741] = 'h000002e5; 	    data_ram[  742] = 'h000002e6; 	    data_ram[  743] = 'h000002e7; 	
    data_ram[  744] = 'h000002e8; 	    data_ram[  745] = 'h000002e9; 	    data_ram[  746] = 'h000002ea; 	    data_ram[  747] = 'h000002eb; 	    data_ram[  748] = 'h000002ec; 	    data_ram[  749] = 'h000002ed; 	    data_ram[  750] = 'h000002ee; 	    data_ram[  751] = 'h000002ef; 	
    data_ram[  752] = 'h000002f0; 	    data_ram[  753] = 'h000002f1; 	    data_ram[  754] = 'h000002f2; 	    data_ram[  755] = 'h000002f3; 	    data_ram[  756] = 'h000002f4; 	    data_ram[  757] = 'h000002f5; 	    data_ram[  758] = 'h000002f6; 	    data_ram[  759] = 'h000002f7; 	
    data_ram[  760] = 'h000002f8; 	    data_ram[  761] = 'h000002f9; 	    data_ram[  762] = 'h000002fa; 	    data_ram[  763] = 'h000002fb; 	    data_ram[  764] = 'h000002fc; 	    data_ram[  765] = 'h000002fd; 	    data_ram[  766] = 'h000002fe; 	    data_ram[  767] = 'h000002ff; 	
    data_ram[  768] = 'h00000300; 	    data_ram[  769] = 'h00000301; 	    data_ram[  770] = 'h00000302; 	    data_ram[  771] = 'h00000303; 	    data_ram[  772] = 'h00000304; 	    data_ram[  773] = 'h00000305; 	    data_ram[  774] = 'h00000306; 	    data_ram[  775] = 'h00000307; 	
    data_ram[  776] = 'h00000308; 	    data_ram[  777] = 'h00000309; 	    data_ram[  778] = 'h0000030a; 	    data_ram[  779] = 'h0000030b; 	    data_ram[  780] = 'h0000030c; 	    data_ram[  781] = 'h0000030d; 	    data_ram[  782] = 'h0000030e; 	    data_ram[  783] = 'h0000030f; 	
    data_ram[  784] = 'h00000310; 	    data_ram[  785] = 'h00000311; 	    data_ram[  786] = 'h00000312; 	    data_ram[  787] = 'h00000313; 	    data_ram[  788] = 'h00000314; 	    data_ram[  789] = 'h00000315; 	    data_ram[  790] = 'h00000316; 	    data_ram[  791] = 'h00000317; 	
    data_ram[  792] = 'h00000318; 	    data_ram[  793] = 'h00000319; 	    data_ram[  794] = 'h0000031a; 	    data_ram[  795] = 'h0000031b; 	    data_ram[  796] = 'h0000031c; 	    data_ram[  797] = 'h0000031d; 	    data_ram[  798] = 'h0000031e; 	    data_ram[  799] = 'h0000031f; 	
    data_ram[  800] = 'h00000320; 	    data_ram[  801] = 'h00000321; 	    data_ram[  802] = 'h00000322; 	    data_ram[  803] = 'h00000323; 	    data_ram[  804] = 'h00000324; 	    data_ram[  805] = 'h00000325; 	    data_ram[  806] = 'h00000326; 	    data_ram[  807] = 'h00000327; 	
    data_ram[  808] = 'h00000328; 	    data_ram[  809] = 'h00000329; 	    data_ram[  810] = 'h0000032a; 	    data_ram[  811] = 'h0000032b; 	    data_ram[  812] = 'h0000032c; 	    data_ram[  813] = 'h0000032d; 	    data_ram[  814] = 'h0000032e; 	    data_ram[  815] = 'h0000032f; 	
    data_ram[  816] = 'h00000330; 	    data_ram[  817] = 'h00000331; 	    data_ram[  818] = 'h00000332; 	    data_ram[  819] = 'h00000333; 	    data_ram[  820] = 'h00000334; 	    data_ram[  821] = 'h00000335; 	    data_ram[  822] = 'h00000336; 	    data_ram[  823] = 'h00000337; 	
    data_ram[  824] = 'h00000338; 	    data_ram[  825] = 'h00000339; 	    data_ram[  826] = 'h0000033a; 	    data_ram[  827] = 'h0000033b; 	    data_ram[  828] = 'h0000033c; 	    data_ram[  829] = 'h0000033d; 	    data_ram[  830] = 'h0000033e; 	    data_ram[  831] = 'h0000033f; 	
    data_ram[  832] = 'h00000340; 	    data_ram[  833] = 'h00000341; 	    data_ram[  834] = 'h00000342; 	    data_ram[  835] = 'h00000343; 	    data_ram[  836] = 'h00000344; 	    data_ram[  837] = 'h00000345; 	    data_ram[  838] = 'h00000346; 	    data_ram[  839] = 'h00000347; 	
    data_ram[  840] = 'h00000348; 	    data_ram[  841] = 'h00000349; 	    data_ram[  842] = 'h0000034a; 	    data_ram[  843] = 'h0000034b; 	    data_ram[  844] = 'h0000034c; 	    data_ram[  845] = 'h0000034d; 	    data_ram[  846] = 'h0000034e; 	    data_ram[  847] = 'h0000034f; 	
    data_ram[  848] = 'h00000350; 	    data_ram[  849] = 'h00000351; 	    data_ram[  850] = 'h00000352; 	    data_ram[  851] = 'h00000353; 	    data_ram[  852] = 'h00000354; 	    data_ram[  853] = 'h00000355; 	    data_ram[  854] = 'h00000356; 	    data_ram[  855] = 'h00000357; 	
    data_ram[  856] = 'h00000358; 	    data_ram[  857] = 'h00000359; 	    data_ram[  858] = 'h0000035a; 	    data_ram[  859] = 'h0000035b; 	    data_ram[  860] = 'h0000035c; 	    data_ram[  861] = 'h0000035d; 	    data_ram[  862] = 'h0000035e; 	    data_ram[  863] = 'h0000035f; 	
    data_ram[  864] = 'h00000360; 	    data_ram[  865] = 'h00000361; 	    data_ram[  866] = 'h00000362; 	    data_ram[  867] = 'h00000363; 	    data_ram[  868] = 'h00000364; 	    data_ram[  869] = 'h00000365; 	    data_ram[  870] = 'h00000366; 	    data_ram[  871] = 'h00000367; 	
    data_ram[  872] = 'h00000368; 	    data_ram[  873] = 'h00000369; 	    data_ram[  874] = 'h0000036a; 	    data_ram[  875] = 'h0000036b; 	    data_ram[  876] = 'h0000036c; 	    data_ram[  877] = 'h0000036d; 	    data_ram[  878] = 'h0000036e; 	    data_ram[  879] = 'h0000036f; 	
    data_ram[  880] = 'h00000370; 	    data_ram[  881] = 'h00000371; 	    data_ram[  882] = 'h00000372; 	    data_ram[  883] = 'h00000373; 	    data_ram[  884] = 'h00000374; 	    data_ram[  885] = 'h00000375; 	    data_ram[  886] = 'h00000376; 	    data_ram[  887] = 'h00000377; 	
    data_ram[  888] = 'h00000378; 	    data_ram[  889] = 'h00000379; 	    data_ram[  890] = 'h0000037a; 	    data_ram[  891] = 'h0000037b; 	    data_ram[  892] = 'h0000037c; 	    data_ram[  893] = 'h0000037d; 	    data_ram[  894] = 'h0000037e; 	    data_ram[  895] = 'h0000037f; 	
    data_ram[  896] = 'h00000380; 	    data_ram[  897] = 'h00000381; 	    data_ram[  898] = 'h00000382; 	    data_ram[  899] = 'h00000383; 	    data_ram[  900] = 'h00000384; 	    data_ram[  901] = 'h00000385; 	    data_ram[  902] = 'h00000386; 	    data_ram[  903] = 'h00000387; 	
    data_ram[  904] = 'h00000388; 	    data_ram[  905] = 'h00000389; 	    data_ram[  906] = 'h0000038a; 	    data_ram[  907] = 'h0000038b; 	    data_ram[  908] = 'h0000038c; 	    data_ram[  909] = 'h0000038d; 	    data_ram[  910] = 'h0000038e; 	    data_ram[  911] = 'h0000038f; 	
    data_ram[  912] = 'h00000390; 	    data_ram[  913] = 'h00000391; 	    data_ram[  914] = 'h00000392; 	    data_ram[  915] = 'h00000393; 	    data_ram[  916] = 'h00000394; 	    data_ram[  917] = 'h00000395; 	    data_ram[  918] = 'h00000396; 	    data_ram[  919] = 'h00000397; 	
    data_ram[  920] = 'h00000398; 	    data_ram[  921] = 'h00000399; 	    data_ram[  922] = 'h0000039a; 	    data_ram[  923] = 'h0000039b; 	    data_ram[  924] = 'h0000039c; 	    data_ram[  925] = 'h0000039d; 	    data_ram[  926] = 'h0000039e; 	    data_ram[  927] = 'h0000039f; 	
    data_ram[  928] = 'h000003a0; 	    data_ram[  929] = 'h000003a1; 	    data_ram[  930] = 'h000003a2; 	    data_ram[  931] = 'h000003a3; 	    data_ram[  932] = 'h000003a4; 	    data_ram[  933] = 'h000003a5; 	    data_ram[  934] = 'h000003a6; 	    data_ram[  935] = 'h000003a7; 	
    data_ram[  936] = 'h000003a8; 	    data_ram[  937] = 'h000003a9; 	    data_ram[  938] = 'h000003aa; 	    data_ram[  939] = 'h000003ab; 	    data_ram[  940] = 'h000003ac; 	    data_ram[  941] = 'h000003ad; 	    data_ram[  942] = 'h000003ae; 	    data_ram[  943] = 'h000003af; 	
    data_ram[  944] = 'h000003b0; 	    data_ram[  945] = 'h000003b1; 	    data_ram[  946] = 'h000003b2; 	    data_ram[  947] = 'h000003b3; 	    data_ram[  948] = 'h000003b4; 	    data_ram[  949] = 'h000003b5; 	    data_ram[  950] = 'h000003b6; 	    data_ram[  951] = 'h000003b7; 	
    data_ram[  952] = 'h000003b8; 	    data_ram[  953] = 'h000003b9; 	    data_ram[  954] = 'h000003ba; 	    data_ram[  955] = 'h000003bb; 	    data_ram[  956] = 'h000003bc; 	    data_ram[  957] = 'h000003bd; 	    data_ram[  958] = 'h000003be; 	    data_ram[  959] = 'h000003bf; 	
    data_ram[  960] = 'h000003c0; 	    data_ram[  961] = 'h000003c1; 	    data_ram[  962] = 'h000003c2; 	    data_ram[  963] = 'h000003c3; 	    data_ram[  964] = 'h000003c4; 	    data_ram[  965] = 'h000003c5; 	    data_ram[  966] = 'h000003c6; 	    data_ram[  967] = 'h000003c7; 	
    data_ram[  968] = 'h000003c8; 	    data_ram[  969] = 'h000003c9; 	    data_ram[  970] = 'h000003ca; 	    data_ram[  971] = 'h000003cb; 	    data_ram[  972] = 'h000003cc; 	    data_ram[  973] = 'h000003cd; 	    data_ram[  974] = 'h000003ce; 	    data_ram[  975] = 'h000003cf; 	
    data_ram[  976] = 'h000003d0; 	    data_ram[  977] = 'h000003d1; 	    data_ram[  978] = 'h000003d2; 	    data_ram[  979] = 'h000003d3; 	    data_ram[  980] = 'h000003d4; 	    data_ram[  981] = 'h000003d5; 	    data_ram[  982] = 'h000003d6; 	    data_ram[  983] = 'h000003d7; 	
    data_ram[  984] = 'h000003d8; 	    data_ram[  985] = 'h000003d9; 	    data_ram[  986] = 'h000003da; 	    data_ram[  987] = 'h000003db; 	    data_ram[  988] = 'h000003dc; 	    data_ram[  989] = 'h000003dd; 	    data_ram[  990] = 'h000003de; 	    data_ram[  991] = 'h000003df; 	
    data_ram[  992] = 'h000003e0; 	    data_ram[  993] = 'h000003e1; 	    data_ram[  994] = 'h000003e2; 	    data_ram[  995] = 'h000003e3; 	    data_ram[  996] = 'h000003e4; 	    data_ram[  997] = 'h000003e5; 	    data_ram[  998] = 'h000003e6; 	    data_ram[  999] = 'h000003e7; 	
    data_ram[ 1000] = 'h000003e8; 	    data_ram[ 1001] = 'h000003e9; 	    data_ram[ 1002] = 'h000003ea; 	    data_ram[ 1003] = 'h000003eb; 	    data_ram[ 1004] = 'h000003ec; 	    data_ram[ 1005] = 'h000003ed; 	    data_ram[ 1006] = 'h000003ee; 	    data_ram[ 1007] = 'h000003ef; 	
    data_ram[ 1008] = 'h000003f0; 	    data_ram[ 1009] = 'h000003f1; 	    data_ram[ 1010] = 'h000003f2; 	    data_ram[ 1011] = 'h000003f3; 	    data_ram[ 1012] = 'h000003f4; 	    data_ram[ 1013] = 'h000003f5; 	    data_ram[ 1014] = 'h000003f6; 	    data_ram[ 1015] = 'h000003f7; 	
    data_ram[ 1016] = 'h000003f8; 	    data_ram[ 1017] = 'h000003f9; 	    data_ram[ 1018] = 'h000003fa; 	    data_ram[ 1019] = 'h000003fb; 	    data_ram[ 1020] = 'h000003fc; 	    data_ram[ 1021] = 'h000003fd; 	    data_ram[ 1022] = 'h000003fe; 	    data_ram[ 1023] = 'h000003ff; 	

end
initial begin
    i_addr_rom[    0] = 'h000002b4; 	    d_addr_rom[    0] = 'h000008ec; 	    wdata_rom[    0] = 'hb0692813; 	    wvalid_rom[    0] = 0; 
    i_addr_rom[    1] = 'h000004d4; 	    d_addr_rom[    1] = 'h00000c34; 	    wdata_rom[    1] = 'h72f0f6fd; 	    wvalid_rom[    1] = 0; 
    i_addr_rom[    2] = 'h000007f8; 	    d_addr_rom[    2] = 'h000009a4; 	    wdata_rom[    2] = 'h2e49ddf3; 	    wvalid_rom[    2] = 0; 
    i_addr_rom[    3] = 'h0000039c; 	    d_addr_rom[    3] = 'h00000e38; 	    wdata_rom[    3] = 'hf55080c7; 	    wvalid_rom[    3] = 0; 
    i_addr_rom[    4] = 'h00000574; 	    d_addr_rom[    4] = 'h00000e2c; 	    wdata_rom[    4] = 'h1dbcb8e8; 	    wvalid_rom[    4] = 1; 
    i_addr_rom[    5] = 'h00000294; 	    d_addr_rom[    5] = 'h00000ce4; 	    wdata_rom[    5] = 'h8307ee13; 	    wvalid_rom[    5] = 1; 
    i_addr_rom[    6] = 'h0000001c; 	    d_addr_rom[    6] = 'h00000820; 	    wdata_rom[    6] = 'hc98db285; 	    wvalid_rom[    6] = 1; 
    i_addr_rom[    7] = 'h00000700; 	    d_addr_rom[    7] = 'h00000c24; 	    wdata_rom[    7] = 'h49daea64; 	    wvalid_rom[    7] = 1; 
    i_addr_rom[    8] = 'h00000074; 	    d_addr_rom[    8] = 'h00000ef8; 	    wdata_rom[    8] = 'h7b163d8e; 	    wvalid_rom[    8] = 0; 
    i_addr_rom[    9] = 'h00000378; 	    d_addr_rom[    9] = 'h000008b0; 	    wdata_rom[    9] = 'h2c016628; 	    wvalid_rom[    9] = 1; 
    i_addr_rom[   10] = 'h000004a0; 	    d_addr_rom[   10] = 'h00000cec; 	    wdata_rom[   10] = 'h9e33ea91; 	    wvalid_rom[   10] = 1; 
    i_addr_rom[   11] = 'h000002c8; 	    d_addr_rom[   11] = 'h00000dc0; 	    wdata_rom[   11] = 'h1dad069d; 	    wvalid_rom[   11] = 1; 
    i_addr_rom[   12] = 'h000005bc; 	    d_addr_rom[   12] = 'h00000bc4; 	    wdata_rom[   12] = 'ha7358d48; 	    wvalid_rom[   12] = 0; 
    i_addr_rom[   13] = 'h00000670; 	    d_addr_rom[   13] = 'h00000f3c; 	    wdata_rom[   13] = 'he211602f; 	    wvalid_rom[   13] = 0; 
    i_addr_rom[   14] = 'h000002a4; 	    d_addr_rom[   14] = 'h00000e80; 	    wdata_rom[   14] = 'he2f10719; 	    wvalid_rom[   14] = 0; 
    i_addr_rom[   15] = 'h00000224; 	    d_addr_rom[   15] = 'h00000e60; 	    wdata_rom[   15] = 'h67e28e06; 	    wvalid_rom[   15] = 0; 
    i_addr_rom[   16] = 'h00000634; 	    d_addr_rom[   16] = 'h00000d4c; 	    wdata_rom[   16] = 'h4741ab9f; 	    wvalid_rom[   16] = 0; 
    i_addr_rom[   17] = 'h0000052c; 	    d_addr_rom[   17] = 'h00000e50; 	    wdata_rom[   17] = 'h67f7b708; 	    wvalid_rom[   17] = 1; 
    i_addr_rom[   18] = 'h0000077c; 	    d_addr_rom[   18] = 'h00000d14; 	    wdata_rom[   18] = 'hdf0e552d; 	    wvalid_rom[   18] = 1; 
    i_addr_rom[   19] = 'h00000708; 	    d_addr_rom[   19] = 'h00000a50; 	    wdata_rom[   19] = 'h0753e227; 	    wvalid_rom[   19] = 0; 
    i_addr_rom[   20] = 'h00000164; 	    d_addr_rom[   20] = 'h000009f4; 	    wdata_rom[   20] = 'h6daa49b9; 	    wvalid_rom[   20] = 0; 
    i_addr_rom[   21] = 'h000001b0; 	    d_addr_rom[   21] = 'h00000c00; 	    wdata_rom[   21] = 'h869ec70d; 	    wvalid_rom[   21] = 0; 
    i_addr_rom[   22] = 'h000002b8; 	    d_addr_rom[   22] = 'h00000b48; 	    wdata_rom[   22] = 'h959fc47b; 	    wvalid_rom[   22] = 0; 
    i_addr_rom[   23] = 'h0000015c; 	    d_addr_rom[   23] = 'h00000c54; 	    wdata_rom[   23] = 'h9a1807cc; 	    wvalid_rom[   23] = 1; 
    i_addr_rom[   24] = 'h000000e4; 	    d_addr_rom[   24] = 'h00000cf4; 	    wdata_rom[   24] = 'h8852b9fa; 	    wvalid_rom[   24] = 1; 
    i_addr_rom[   25] = 'h000003b0; 	    d_addr_rom[   25] = 'h0000099c; 	    wdata_rom[   25] = 'hdfec1e9d; 	    wvalid_rom[   25] = 1; 
    i_addr_rom[   26] = 'h00000310; 	    d_addr_rom[   26] = 'h000008c8; 	    wdata_rom[   26] = 'h5cf71411; 	    wvalid_rom[   26] = 1; 
    i_addr_rom[   27] = 'h000006a4; 	    d_addr_rom[   27] = 'h00000c6c; 	    wdata_rom[   27] = 'hf0a45954; 	    wvalid_rom[   27] = 0; 
    i_addr_rom[   28] = 'h00000548; 	    d_addr_rom[   28] = 'h00000a0c; 	    wdata_rom[   28] = 'h3975f64f; 	    wvalid_rom[   28] = 0; 
    i_addr_rom[   29] = 'h000002a8; 	    d_addr_rom[   29] = 'h00000bfc; 	    wdata_rom[   29] = 'h04f069b9; 	    wvalid_rom[   29] = 1; 
    i_addr_rom[   30] = 'h000002ac; 	    d_addr_rom[   30] = 'h00000e60; 	    wdata_rom[   30] = 'h7ba891e4; 	    wvalid_rom[   30] = 1; 
    i_addr_rom[   31] = 'h00000750; 	    d_addr_rom[   31] = 'h00000f6c; 	    wdata_rom[   31] = 'h6ef28e83; 	    wvalid_rom[   31] = 1; 
    i_addr_rom[   32] = 'h00000714; 	    d_addr_rom[   32] = 'h00000a38; 	    wdata_rom[   32] = 'h85e5db9c; 	    wvalid_rom[   32] = 0; 
    i_addr_rom[   33] = 'h00000330; 	    d_addr_rom[   33] = 'h00000e34; 	    wdata_rom[   33] = 'hd32438ac; 	    wvalid_rom[   33] = 1; 
    i_addr_rom[   34] = 'h000003c8; 	    d_addr_rom[   34] = 'h00000f04; 	    wdata_rom[   34] = 'h96e0b9dd; 	    wvalid_rom[   34] = 1; 
    i_addr_rom[   35] = 'h00000610; 	    d_addr_rom[   35] = 'h00000d8c; 	    wdata_rom[   35] = 'h2693e698; 	    wvalid_rom[   35] = 0; 
    i_addr_rom[   36] = 'h0000074c; 	    d_addr_rom[   36] = 'h00000d38; 	    wdata_rom[   36] = 'hc92b9c1c; 	    wvalid_rom[   36] = 0; 
    i_addr_rom[   37] = 'h00000598; 	    d_addr_rom[   37] = 'h00000dd4; 	    wdata_rom[   37] = 'hc817eb20; 	    wvalid_rom[   37] = 1; 
    i_addr_rom[   38] = 'h000007e8; 	    d_addr_rom[   38] = 'h00000994; 	    wdata_rom[   38] = 'h94a577dd; 	    wvalid_rom[   38] = 0; 
    i_addr_rom[   39] = 'h00000148; 	    d_addr_rom[   39] = 'h00000afc; 	    wdata_rom[   39] = 'h3e2f0c47; 	    wvalid_rom[   39] = 1; 
    i_addr_rom[   40] = 'h00000108; 	    d_addr_rom[   40] = 'h00000934; 	    wdata_rom[   40] = 'h31e6b9c3; 	    wvalid_rom[   40] = 0; 
    i_addr_rom[   41] = 'h000005b8; 	    d_addr_rom[   41] = 'h000008ec; 	    wdata_rom[   41] = 'hb69e041a; 	    wvalid_rom[   41] = 1; 
    i_addr_rom[   42] = 'h000000a4; 	    d_addr_rom[   42] = 'h00000b30; 	    wdata_rom[   42] = 'he1735815; 	    wvalid_rom[   42] = 1; 
    i_addr_rom[   43] = 'h000001e4; 	    d_addr_rom[   43] = 'h00000860; 	    wdata_rom[   43] = 'hdf8eee56; 	    wvalid_rom[   43] = 0; 
    i_addr_rom[   44] = 'h000007c4; 	    d_addr_rom[   44] = 'h00000834; 	    wdata_rom[   44] = 'he0f4fbfc; 	    wvalid_rom[   44] = 1; 
    i_addr_rom[   45] = 'h00000134; 	    d_addr_rom[   45] = 'h00000e20; 	    wdata_rom[   45] = 'h13b45062; 	    wvalid_rom[   45] = 0; 
    i_addr_rom[   46] = 'h0000071c; 	    d_addr_rom[   46] = 'h00000d70; 	    wdata_rom[   46] = 'h58a1065f; 	    wvalid_rom[   46] = 1; 
    i_addr_rom[   47] = 'h00000240; 	    d_addr_rom[   47] = 'h00000d80; 	    wdata_rom[   47] = 'hede62fcb; 	    wvalid_rom[   47] = 1; 
    i_addr_rom[   48] = 'h000002f0; 	    d_addr_rom[   48] = 'h00000eb4; 	    wdata_rom[   48] = 'h7edd89e8; 	    wvalid_rom[   48] = 1; 
    i_addr_rom[   49] = 'h0000055c; 	    d_addr_rom[   49] = 'h00000b58; 	    wdata_rom[   49] = 'h4bbd0ea7; 	    wvalid_rom[   49] = 0; 
    i_addr_rom[   50] = 'h00000474; 	    d_addr_rom[   50] = 'h00000fec; 	    wdata_rom[   50] = 'h439fdb55; 	    wvalid_rom[   50] = 1; 
    i_addr_rom[   51] = 'h00000104; 	    d_addr_rom[   51] = 'h00000d00; 	    wdata_rom[   51] = 'hff046c90; 	    wvalid_rom[   51] = 0; 
    i_addr_rom[   52] = 'h0000037c; 	    d_addr_rom[   52] = 'h000009d8; 	    wdata_rom[   52] = 'h5d0018e3; 	    wvalid_rom[   52] = 1; 
    i_addr_rom[   53] = 'h0000068c; 	    d_addr_rom[   53] = 'h00000870; 	    wdata_rom[   53] = 'h1d28a8db; 	    wvalid_rom[   53] = 0; 
    i_addr_rom[   54] = 'h00000688; 	    d_addr_rom[   54] = 'h00000a28; 	    wdata_rom[   54] = 'h8d70b05b; 	    wvalid_rom[   54] = 1; 
    i_addr_rom[   55] = 'h00000658; 	    d_addr_rom[   55] = 'h00000eec; 	    wdata_rom[   55] = 'h6c99a1cb; 	    wvalid_rom[   55] = 0; 
    i_addr_rom[   56] = 'h0000017c; 	    d_addr_rom[   56] = 'h000009a0; 	    wdata_rom[   56] = 'h9cddd433; 	    wvalid_rom[   56] = 0; 
    i_addr_rom[   57] = 'h0000069c; 	    d_addr_rom[   57] = 'h000008d8; 	    wdata_rom[   57] = 'h027b2f3e; 	    wvalid_rom[   57] = 1; 
    i_addr_rom[   58] = 'h00000298; 	    d_addr_rom[   58] = 'h00000e70; 	    wdata_rom[   58] = 'h5fe86bbd; 	    wvalid_rom[   58] = 0; 
    i_addr_rom[   59] = 'h0000021c; 	    d_addr_rom[   59] = 'h00000a98; 	    wdata_rom[   59] = 'ha86d9e8c; 	    wvalid_rom[   59] = 0; 
    i_addr_rom[   60] = 'h0000027c; 	    d_addr_rom[   60] = 'h00000cd0; 	    wdata_rom[   60] = 'hfaa1ce1b; 	    wvalid_rom[   60] = 1; 
    i_addr_rom[   61] = 'h000001bc; 	    d_addr_rom[   61] = 'h00000c3c; 	    wdata_rom[   61] = 'h492c0867; 	    wvalid_rom[   61] = 0; 
    i_addr_rom[   62] = 'h00000180; 	    d_addr_rom[   62] = 'h00000bac; 	    wdata_rom[   62] = 'h40bba9d4; 	    wvalid_rom[   62] = 1; 
    i_addr_rom[   63] = 'h00000418; 	    d_addr_rom[   63] = 'h00000ca0; 	    wdata_rom[   63] = 'hd590eba0; 	    wvalid_rom[   63] = 0; 
    i_addr_rom[   64] = 'h00000410; 	    d_addr_rom[   64] = 'h00000fc8; 	    wdata_rom[   64] = 'h0818e257; 	    wvalid_rom[   64] = 0; 
    i_addr_rom[   65] = 'h00000748; 	    d_addr_rom[   65] = 'h00000bd4; 	    wdata_rom[   65] = 'h32e5692f; 	    wvalid_rom[   65] = 0; 
    i_addr_rom[   66] = 'h00000280; 	    d_addr_rom[   66] = 'h00000d0c; 	    wdata_rom[   66] = 'hea9c9023; 	    wvalid_rom[   66] = 0; 
    i_addr_rom[   67] = 'h00000228; 	    d_addr_rom[   67] = 'h00000dd8; 	    wdata_rom[   67] = 'ha597aea4; 	    wvalid_rom[   67] = 0; 
    i_addr_rom[   68] = 'h00000088; 	    d_addr_rom[   68] = 'h00000a54; 	    wdata_rom[   68] = 'h57442387; 	    wvalid_rom[   68] = 1; 
    i_addr_rom[   69] = 'h00000708; 	    d_addr_rom[   69] = 'h00000dc4; 	    wdata_rom[   69] = 'h928e9687; 	    wvalid_rom[   69] = 0; 
    i_addr_rom[   70] = 'h000003a0; 	    d_addr_rom[   70] = 'h00000f50; 	    wdata_rom[   70] = 'hb38b97e1; 	    wvalid_rom[   70] = 0; 
    i_addr_rom[   71] = 'h000000e0; 	    d_addr_rom[   71] = 'h00000abc; 	    wdata_rom[   71] = 'h0c58fc95; 	    wvalid_rom[   71] = 0; 
    i_addr_rom[   72] = 'h00000460; 	    d_addr_rom[   72] = 'h00000b68; 	    wdata_rom[   72] = 'hc652d8fb; 	    wvalid_rom[   72] = 1; 
    i_addr_rom[   73] = 'h000005cc; 	    d_addr_rom[   73] = 'h000009b4; 	    wdata_rom[   73] = 'he48d2078; 	    wvalid_rom[   73] = 1; 
    i_addr_rom[   74] = 'h00000654; 	    d_addr_rom[   74] = 'h00000d0c; 	    wdata_rom[   74] = 'hb16c32d3; 	    wvalid_rom[   74] = 1; 
    i_addr_rom[   75] = 'h00000378; 	    d_addr_rom[   75] = 'h00000830; 	    wdata_rom[   75] = 'h5c7a58e7; 	    wvalid_rom[   75] = 0; 
    i_addr_rom[   76] = 'h0000024c; 	    d_addr_rom[   76] = 'h00000d70; 	    wdata_rom[   76] = 'h910a8712; 	    wvalid_rom[   76] = 1; 
    i_addr_rom[   77] = 'h000002ac; 	    d_addr_rom[   77] = 'h00000fdc; 	    wdata_rom[   77] = 'h90d3000c; 	    wvalid_rom[   77] = 0; 
    i_addr_rom[   78] = 'h000005f4; 	    d_addr_rom[   78] = 'h000008fc; 	    wdata_rom[   78] = 'h1ca72eaf; 	    wvalid_rom[   78] = 0; 
    i_addr_rom[   79] = 'h0000020c; 	    d_addr_rom[   79] = 'h00000b50; 	    wdata_rom[   79] = 'h1d09a11b; 	    wvalid_rom[   79] = 0; 
    i_addr_rom[   80] = 'h00000718; 	    d_addr_rom[   80] = 'h000009a0; 	    wdata_rom[   80] = 'h87bab5bc; 	    wvalid_rom[   80] = 0; 
    i_addr_rom[   81] = 'h00000220; 	    d_addr_rom[   81] = 'h00000d34; 	    wdata_rom[   81] = 'h79d805b9; 	    wvalid_rom[   81] = 0; 
    i_addr_rom[   82] = 'h0000056c; 	    d_addr_rom[   82] = 'h00000de8; 	    wdata_rom[   82] = 'h460bef80; 	    wvalid_rom[   82] = 1; 
    i_addr_rom[   83] = 'h000006fc; 	    d_addr_rom[   83] = 'h00000d14; 	    wdata_rom[   83] = 'hd369d116; 	    wvalid_rom[   83] = 1; 
    i_addr_rom[   84] = 'h000003ec; 	    d_addr_rom[   84] = 'h00000fe4; 	    wdata_rom[   84] = 'h82babbd9; 	    wvalid_rom[   84] = 1; 
    i_addr_rom[   85] = 'h00000018; 	    d_addr_rom[   85] = 'h00000878; 	    wdata_rom[   85] = 'h385a248f; 	    wvalid_rom[   85] = 0; 
    i_addr_rom[   86] = 'h00000598; 	    d_addr_rom[   86] = 'h00000808; 	    wdata_rom[   86] = 'h7a722eb6; 	    wvalid_rom[   86] = 1; 
    i_addr_rom[   87] = 'h00000664; 	    d_addr_rom[   87] = 'h00000ac8; 	    wdata_rom[   87] = 'hb496456f; 	    wvalid_rom[   87] = 1; 
    i_addr_rom[   88] = 'h000004d4; 	    d_addr_rom[   88] = 'h00000a74; 	    wdata_rom[   88] = 'hefc0dfb7; 	    wvalid_rom[   88] = 0; 
    i_addr_rom[   89] = 'h00000270; 	    d_addr_rom[   89] = 'h00000eb8; 	    wdata_rom[   89] = 'h249d7a2b; 	    wvalid_rom[   89] = 0; 
    i_addr_rom[   90] = 'h00000690; 	    d_addr_rom[   90] = 'h000009b0; 	    wdata_rom[   90] = 'h56d60792; 	    wvalid_rom[   90] = 1; 
    i_addr_rom[   91] = 'h000000d8; 	    d_addr_rom[   91] = 'h00000958; 	    wdata_rom[   91] = 'h4594876a; 	    wvalid_rom[   91] = 0; 
    i_addr_rom[   92] = 'h0000022c; 	    d_addr_rom[   92] = 'h00000d70; 	    wdata_rom[   92] = 'hb2d2ac10; 	    wvalid_rom[   92] = 0; 
    i_addr_rom[   93] = 'h000007e8; 	    d_addr_rom[   93] = 'h00000990; 	    wdata_rom[   93] = 'h626e5ce9; 	    wvalid_rom[   93] = 1; 
    i_addr_rom[   94] = 'h0000006c; 	    d_addr_rom[   94] = 'h00000da0; 	    wdata_rom[   94] = 'h7942eca1; 	    wvalid_rom[   94] = 0; 
    i_addr_rom[   95] = 'h00000318; 	    d_addr_rom[   95] = 'h00000acc; 	    wdata_rom[   95] = 'h2b6542d3; 	    wvalid_rom[   95] = 1; 
    i_addr_rom[   96] = 'h00000794; 	    d_addr_rom[   96] = 'h00000860; 	    wdata_rom[   96] = 'h4103a792; 	    wvalid_rom[   96] = 0; 
    i_addr_rom[   97] = 'h000003f4; 	    d_addr_rom[   97] = 'h00000adc; 	    wdata_rom[   97] = 'h887ca6df; 	    wvalid_rom[   97] = 0; 
    i_addr_rom[   98] = 'h000000c8; 	    d_addr_rom[   98] = 'h00000d50; 	    wdata_rom[   98] = 'hde796b8e; 	    wvalid_rom[   98] = 1; 
    i_addr_rom[   99] = 'h000004b8; 	    d_addr_rom[   99] = 'h00000918; 	    wdata_rom[   99] = 'h16b98ff2; 	    wvalid_rom[   99] = 0; 
    i_addr_rom[  100] = 'h000002d0; 	    d_addr_rom[  100] = 'h00000e5c; 	    wdata_rom[  100] = 'h1409852d; 	    wvalid_rom[  100] = 1; 
    i_addr_rom[  101] = 'h000003c0; 	    d_addr_rom[  101] = 'h00000f24; 	    wdata_rom[  101] = 'hcecd7e4d; 	    wvalid_rom[  101] = 1; 
    i_addr_rom[  102] = 'h00000458; 	    d_addr_rom[  102] = 'h000008d4; 	    wdata_rom[  102] = 'h2fbf4a87; 	    wvalid_rom[  102] = 0; 
    i_addr_rom[  103] = 'h00000238; 	    d_addr_rom[  103] = 'h000009ac; 	    wdata_rom[  103] = 'h1ddf08de; 	    wvalid_rom[  103] = 1; 
    i_addr_rom[  104] = 'h000004ec; 	    d_addr_rom[  104] = 'h00000884; 	    wdata_rom[  104] = 'h5380ae9e; 	    wvalid_rom[  104] = 0; 
    i_addr_rom[  105] = 'h0000071c; 	    d_addr_rom[  105] = 'h00000ab4; 	    wdata_rom[  105] = 'h3cd8d32d; 	    wvalid_rom[  105] = 0; 
    i_addr_rom[  106] = 'h000006d8; 	    d_addr_rom[  106] = 'h000009f0; 	    wdata_rom[  106] = 'h40056275; 	    wvalid_rom[  106] = 0; 
    i_addr_rom[  107] = 'h0000023c; 	    d_addr_rom[  107] = 'h00000a10; 	    wdata_rom[  107] = 'he3380a6c; 	    wvalid_rom[  107] = 0; 
    i_addr_rom[  108] = 'h00000514; 	    d_addr_rom[  108] = 'h00000c74; 	    wdata_rom[  108] = 'hcf4188c5; 	    wvalid_rom[  108] = 0; 
    i_addr_rom[  109] = 'h0000079c; 	    d_addr_rom[  109] = 'h00000ddc; 	    wdata_rom[  109] = 'h48386f41; 	    wvalid_rom[  109] = 1; 
    i_addr_rom[  110] = 'h0000001c; 	    d_addr_rom[  110] = 'h00000f44; 	    wdata_rom[  110] = 'h68bdb77d; 	    wvalid_rom[  110] = 0; 
    i_addr_rom[  111] = 'h000000e8; 	    d_addr_rom[  111] = 'h00000ab0; 	    wdata_rom[  111] = 'hd481428c; 	    wvalid_rom[  111] = 1; 
    i_addr_rom[  112] = 'h000002d4; 	    d_addr_rom[  112] = 'h00000b04; 	    wdata_rom[  112] = 'hb27f4e9c; 	    wvalid_rom[  112] = 0; 
    i_addr_rom[  113] = 'h00000484; 	    d_addr_rom[  113] = 'h00000e70; 	    wdata_rom[  113] = 'h19c00014; 	    wvalid_rom[  113] = 0; 
    i_addr_rom[  114] = 'h00000014; 	    d_addr_rom[  114] = 'h00000eb4; 	    wdata_rom[  114] = 'hb4fbdb7b; 	    wvalid_rom[  114] = 1; 
    i_addr_rom[  115] = 'h00000084; 	    d_addr_rom[  115] = 'h00000aec; 	    wdata_rom[  115] = 'h68cc5975; 	    wvalid_rom[  115] = 1; 
    i_addr_rom[  116] = 'h000004c0; 	    d_addr_rom[  116] = 'h00000e78; 	    wdata_rom[  116] = 'h8e755d7c; 	    wvalid_rom[  116] = 0; 
    i_addr_rom[  117] = 'h00000258; 	    d_addr_rom[  117] = 'h00000d78; 	    wdata_rom[  117] = 'h5864aef4; 	    wvalid_rom[  117] = 1; 
    i_addr_rom[  118] = 'h0000022c; 	    d_addr_rom[  118] = 'h00000e5c; 	    wdata_rom[  118] = 'hcebbb038; 	    wvalid_rom[  118] = 1; 
    i_addr_rom[  119] = 'h00000404; 	    d_addr_rom[  119] = 'h00000908; 	    wdata_rom[  119] = 'h2cf49c61; 	    wvalid_rom[  119] = 1; 
    i_addr_rom[  120] = 'h00000678; 	    d_addr_rom[  120] = 'h00000c64; 	    wdata_rom[  120] = 'h9eaf7ef9; 	    wvalid_rom[  120] = 0; 
    i_addr_rom[  121] = 'h00000364; 	    d_addr_rom[  121] = 'h00000c80; 	    wdata_rom[  121] = 'hb13c1e3b; 	    wvalid_rom[  121] = 1; 
    i_addr_rom[  122] = 'h000001fc; 	    d_addr_rom[  122] = 'h000009d4; 	    wdata_rom[  122] = 'he47ce669; 	    wvalid_rom[  122] = 0; 
    i_addr_rom[  123] = 'h000007c0; 	    d_addr_rom[  123] = 'h00000bc4; 	    wdata_rom[  123] = 'hf1a1bb19; 	    wvalid_rom[  123] = 0; 
    i_addr_rom[  124] = 'h00000390; 	    d_addr_rom[  124] = 'h00000f64; 	    wdata_rom[  124] = 'h5f00c5de; 	    wvalid_rom[  124] = 0; 
    i_addr_rom[  125] = 'h0000065c; 	    d_addr_rom[  125] = 'h00000870; 	    wdata_rom[  125] = 'hb4059d98; 	    wvalid_rom[  125] = 1; 
    i_addr_rom[  126] = 'h0000030c; 	    d_addr_rom[  126] = 'h0000084c; 	    wdata_rom[  126] = 'h22f33bbb; 	    wvalid_rom[  126] = 0; 
    i_addr_rom[  127] = 'h00000764; 	    d_addr_rom[  127] = 'h00000a24; 	    wdata_rom[  127] = 'h5ece1d18; 	    wvalid_rom[  127] = 0; 
    i_addr_rom[  128] = 'h00000304; 	    d_addr_rom[  128] = 'h0000093c; 	    wdata_rom[  128] = 'h2e804494; 	    wvalid_rom[  128] = 0; 
    i_addr_rom[  129] = 'h000004ac; 	    d_addr_rom[  129] = 'h00000e64; 	    wdata_rom[  129] = 'hd4426356; 	    wvalid_rom[  129] = 1; 
    i_addr_rom[  130] = 'h00000214; 	    d_addr_rom[  130] = 'h0000087c; 	    wdata_rom[  130] = 'h778adfaa; 	    wvalid_rom[  130] = 0; 
    i_addr_rom[  131] = 'h0000065c; 	    d_addr_rom[  131] = 'h00000d84; 	    wdata_rom[  131] = 'he0e2b5bf; 	    wvalid_rom[  131] = 0; 
    i_addr_rom[  132] = 'h00000040; 	    d_addr_rom[  132] = 'h00000e40; 	    wdata_rom[  132] = 'hccfd07a4; 	    wvalid_rom[  132] = 1; 
    i_addr_rom[  133] = 'h000000c8; 	    d_addr_rom[  133] = 'h00000be4; 	    wdata_rom[  133] = 'h2a260d62; 	    wvalid_rom[  133] = 0; 
    i_addr_rom[  134] = 'h000005ac; 	    d_addr_rom[  134] = 'h00000970; 	    wdata_rom[  134] = 'hc78208d3; 	    wvalid_rom[  134] = 1; 
    i_addr_rom[  135] = 'h00000728; 	    d_addr_rom[  135] = 'h00000a8c; 	    wdata_rom[  135] = 'h7f2deae7; 	    wvalid_rom[  135] = 0; 
    i_addr_rom[  136] = 'h00000690; 	    d_addr_rom[  136] = 'h00000a18; 	    wdata_rom[  136] = 'h58dd3fec; 	    wvalid_rom[  136] = 1; 
    i_addr_rom[  137] = 'h000005b4; 	    d_addr_rom[  137] = 'h00000b64; 	    wdata_rom[  137] = 'h80a66788; 	    wvalid_rom[  137] = 0; 
    i_addr_rom[  138] = 'h00000148; 	    d_addr_rom[  138] = 'h000008b0; 	    wdata_rom[  138] = 'h2d033e30; 	    wvalid_rom[  138] = 0; 
    i_addr_rom[  139] = 'h00000518; 	    d_addr_rom[  139] = 'h00000ea8; 	    wdata_rom[  139] = 'hbdbfff65; 	    wvalid_rom[  139] = 0; 
    i_addr_rom[  140] = 'h00000440; 	    d_addr_rom[  140] = 'h000009e0; 	    wdata_rom[  140] = 'h18c5febc; 	    wvalid_rom[  140] = 1; 
    i_addr_rom[  141] = 'h000001a4; 	    d_addr_rom[  141] = 'h00000970; 	    wdata_rom[  141] = 'hfd4e31de; 	    wvalid_rom[  141] = 0; 
    i_addr_rom[  142] = 'h000006a4; 	    d_addr_rom[  142] = 'h00000fb0; 	    wdata_rom[  142] = 'h09fcf2a3; 	    wvalid_rom[  142] = 0; 
    i_addr_rom[  143] = 'h0000077c; 	    d_addr_rom[  143] = 'h00000948; 	    wdata_rom[  143] = 'hfd86974b; 	    wvalid_rom[  143] = 0; 
    i_addr_rom[  144] = 'h000000dc; 	    d_addr_rom[  144] = 'h00000844; 	    wdata_rom[  144] = 'hf260bf97; 	    wvalid_rom[  144] = 1; 
    i_addr_rom[  145] = 'h00000144; 	    d_addr_rom[  145] = 'h000009fc; 	    wdata_rom[  145] = 'hea5374d3; 	    wvalid_rom[  145] = 1; 
    i_addr_rom[  146] = 'h000007f0; 	    d_addr_rom[  146] = 'h00000f04; 	    wdata_rom[  146] = 'h971774c2; 	    wvalid_rom[  146] = 0; 
    i_addr_rom[  147] = 'h000005b4; 	    d_addr_rom[  147] = 'h00000d90; 	    wdata_rom[  147] = 'h64a32b8c; 	    wvalid_rom[  147] = 0; 
    i_addr_rom[  148] = 'h0000033c; 	    d_addr_rom[  148] = 'h000009ac; 	    wdata_rom[  148] = 'h0e6198c1; 	    wvalid_rom[  148] = 0; 
    i_addr_rom[  149] = 'h00000090; 	    d_addr_rom[  149] = 'h00000f44; 	    wdata_rom[  149] = 'hff86a389; 	    wvalid_rom[  149] = 1; 
    i_addr_rom[  150] = 'h00000194; 	    d_addr_rom[  150] = 'h00000bd0; 	    wdata_rom[  150] = 'hca2387bd; 	    wvalid_rom[  150] = 0; 
    i_addr_rom[  151] = 'h00000548; 	    d_addr_rom[  151] = 'h00000838; 	    wdata_rom[  151] = 'h3ad948c5; 	    wvalid_rom[  151] = 1; 
    i_addr_rom[  152] = 'h000004cc; 	    d_addr_rom[  152] = 'h00000f84; 	    wdata_rom[  152] = 'h6cafa2df; 	    wvalid_rom[  152] = 0; 
    i_addr_rom[  153] = 'h00000004; 	    d_addr_rom[  153] = 'h00000b20; 	    wdata_rom[  153] = 'hd4185bf0; 	    wvalid_rom[  153] = 0; 
    i_addr_rom[  154] = 'h000005b8; 	    d_addr_rom[  154] = 'h00000da8; 	    wdata_rom[  154] = 'h53dacdf8; 	    wvalid_rom[  154] = 1; 
    i_addr_rom[  155] = 'h00000444; 	    d_addr_rom[  155] = 'h00000d00; 	    wdata_rom[  155] = 'hc518d947; 	    wvalid_rom[  155] = 1; 
    i_addr_rom[  156] = 'h000007b4; 	    d_addr_rom[  156] = 'h000008d0; 	    wdata_rom[  156] = 'h45ec0f13; 	    wvalid_rom[  156] = 0; 
    i_addr_rom[  157] = 'h00000464; 	    d_addr_rom[  157] = 'h00000e8c; 	    wdata_rom[  157] = 'h37368f5f; 	    wvalid_rom[  157] = 0; 
    i_addr_rom[  158] = 'h0000037c; 	    d_addr_rom[  158] = 'h000009bc; 	    wdata_rom[  158] = 'h7102dbfa; 	    wvalid_rom[  158] = 0; 
    i_addr_rom[  159] = 'h00000570; 	    d_addr_rom[  159] = 'h00000f58; 	    wdata_rom[  159] = 'hc7a513e4; 	    wvalid_rom[  159] = 0; 
    i_addr_rom[  160] = 'h00000548; 	    d_addr_rom[  160] = 'h00000c40; 	    wdata_rom[  160] = 'h2e8ac55a; 	    wvalid_rom[  160] = 1; 
    i_addr_rom[  161] = 'h000003b4; 	    d_addr_rom[  161] = 'h00000fdc; 	    wdata_rom[  161] = 'h25b3920b; 	    wvalid_rom[  161] = 1; 
    i_addr_rom[  162] = 'h00000380; 	    d_addr_rom[  162] = 'h00000898; 	    wdata_rom[  162] = 'h93bc8656; 	    wvalid_rom[  162] = 0; 
    i_addr_rom[  163] = 'h00000014; 	    d_addr_rom[  163] = 'h000008e8; 	    wdata_rom[  163] = 'h06d7f2cd; 	    wvalid_rom[  163] = 0; 
    i_addr_rom[  164] = 'h0000009c; 	    d_addr_rom[  164] = 'h00000b6c; 	    wdata_rom[  164] = 'h7e3a958b; 	    wvalid_rom[  164] = 0; 
    i_addr_rom[  165] = 'h000007dc; 	    d_addr_rom[  165] = 'h00000fd8; 	    wdata_rom[  165] = 'hd2d908d0; 	    wvalid_rom[  165] = 1; 
    i_addr_rom[  166] = 'h00000394; 	    d_addr_rom[  166] = 'h00000c04; 	    wdata_rom[  166] = 'h2495ebf7; 	    wvalid_rom[  166] = 1; 
    i_addr_rom[  167] = 'h00000584; 	    d_addr_rom[  167] = 'h00000940; 	    wdata_rom[  167] = 'h1df0370e; 	    wvalid_rom[  167] = 1; 
    i_addr_rom[  168] = 'h000006c4; 	    d_addr_rom[  168] = 'h00000b60; 	    wdata_rom[  168] = 'h554250b8; 	    wvalid_rom[  168] = 0; 
    i_addr_rom[  169] = 'h0000078c; 	    d_addr_rom[  169] = 'h00000ee0; 	    wdata_rom[  169] = 'h46134e21; 	    wvalid_rom[  169] = 1; 
    i_addr_rom[  170] = 'h00000234; 	    d_addr_rom[  170] = 'h00000c50; 	    wdata_rom[  170] = 'hdbbb4ea4; 	    wvalid_rom[  170] = 0; 
    i_addr_rom[  171] = 'h0000036c; 	    d_addr_rom[  171] = 'h00000e90; 	    wdata_rom[  171] = 'h04a27f25; 	    wvalid_rom[  171] = 1; 
    i_addr_rom[  172] = 'h00000144; 	    d_addr_rom[  172] = 'h00000acc; 	    wdata_rom[  172] = 'h85fa3618; 	    wvalid_rom[  172] = 0; 
    i_addr_rom[  173] = 'h00000700; 	    d_addr_rom[  173] = 'h00000b28; 	    wdata_rom[  173] = 'ha274c4f6; 	    wvalid_rom[  173] = 1; 
    i_addr_rom[  174] = 'h000002f0; 	    d_addr_rom[  174] = 'h00000ddc; 	    wdata_rom[  174] = 'haade889c; 	    wvalid_rom[  174] = 0; 
    i_addr_rom[  175] = 'h000004e8; 	    d_addr_rom[  175] = 'h00000f94; 	    wdata_rom[  175] = 'h7faa5578; 	    wvalid_rom[  175] = 1; 
    i_addr_rom[  176] = 'h00000190; 	    d_addr_rom[  176] = 'h00000f54; 	    wdata_rom[  176] = 'h4134e2f0; 	    wvalid_rom[  176] = 1; 
    i_addr_rom[  177] = 'h0000004c; 	    d_addr_rom[  177] = 'h00000a08; 	    wdata_rom[  177] = 'h3613d06f; 	    wvalid_rom[  177] = 1; 
    i_addr_rom[  178] = 'h000002f4; 	    d_addr_rom[  178] = 'h00000978; 	    wdata_rom[  178] = 'h7b240f20; 	    wvalid_rom[  178] = 0; 
    i_addr_rom[  179] = 'h0000052c; 	    d_addr_rom[  179] = 'h00000b28; 	    wdata_rom[  179] = 'h7bc2c916; 	    wvalid_rom[  179] = 1; 
    i_addr_rom[  180] = 'h0000012c; 	    d_addr_rom[  180] = 'h00000858; 	    wdata_rom[  180] = 'h40ad4397; 	    wvalid_rom[  180] = 1; 
    i_addr_rom[  181] = 'h000002b0; 	    d_addr_rom[  181] = 'h0000096c; 	    wdata_rom[  181] = 'hcb042c87; 	    wvalid_rom[  181] = 0; 
    i_addr_rom[  182] = 'h0000079c; 	    d_addr_rom[  182] = 'h00000848; 	    wdata_rom[  182] = 'h331bc675; 	    wvalid_rom[  182] = 0; 
    i_addr_rom[  183] = 'h00000598; 	    d_addr_rom[  183] = 'h00000c18; 	    wdata_rom[  183] = 'hfc1d133e; 	    wvalid_rom[  183] = 1; 
    i_addr_rom[  184] = 'h00000278; 	    d_addr_rom[  184] = 'h000009d4; 	    wdata_rom[  184] = 'h22ade07f; 	    wvalid_rom[  184] = 1; 
    i_addr_rom[  185] = 'h00000058; 	    d_addr_rom[  185] = 'h00000fa8; 	    wdata_rom[  185] = 'h8c27faf1; 	    wvalid_rom[  185] = 0; 
    i_addr_rom[  186] = 'h000001a4; 	    d_addr_rom[  186] = 'h00000830; 	    wdata_rom[  186] = 'h48640243; 	    wvalid_rom[  186] = 0; 
    i_addr_rom[  187] = 'h0000065c; 	    d_addr_rom[  187] = 'h000009f4; 	    wdata_rom[  187] = 'h8811215d; 	    wvalid_rom[  187] = 1; 
    i_addr_rom[  188] = 'h000002f4; 	    d_addr_rom[  188] = 'h00000948; 	    wdata_rom[  188] = 'hb9110d6f; 	    wvalid_rom[  188] = 1; 
    i_addr_rom[  189] = 'h000002a8; 	    d_addr_rom[  189] = 'h00000aac; 	    wdata_rom[  189] = 'h9133e4f6; 	    wvalid_rom[  189] = 0; 
    i_addr_rom[  190] = 'h00000068; 	    d_addr_rom[  190] = 'h00000d70; 	    wdata_rom[  190] = 'ha0c883f6; 	    wvalid_rom[  190] = 1; 
    i_addr_rom[  191] = 'h000000a4; 	    d_addr_rom[  191] = 'h00000b14; 	    wdata_rom[  191] = 'h85a88ab2; 	    wvalid_rom[  191] = 1; 
    i_addr_rom[  192] = 'h00000570; 	    d_addr_rom[  192] = 'h00000b90; 	    wdata_rom[  192] = 'ha54d4eab; 	    wvalid_rom[  192] = 1; 
    i_addr_rom[  193] = 'h0000009c; 	    d_addr_rom[  193] = 'h00000d40; 	    wdata_rom[  193] = 'hd1842f49; 	    wvalid_rom[  193] = 0; 
    i_addr_rom[  194] = 'h0000055c; 	    d_addr_rom[  194] = 'h00000cc0; 	    wdata_rom[  194] = 'h1db8097d; 	    wvalid_rom[  194] = 0; 
    i_addr_rom[  195] = 'h0000026c; 	    d_addr_rom[  195] = 'h00000a04; 	    wdata_rom[  195] = 'h0f5b7341; 	    wvalid_rom[  195] = 0; 
    i_addr_rom[  196] = 'h00000264; 	    d_addr_rom[  196] = 'h00000e6c; 	    wdata_rom[  196] = 'h2b44f98b; 	    wvalid_rom[  196] = 0; 
    i_addr_rom[  197] = 'h00000450; 	    d_addr_rom[  197] = 'h00000bcc; 	    wdata_rom[  197] = 'h141fa03c; 	    wvalid_rom[  197] = 0; 
    i_addr_rom[  198] = 'h0000059c; 	    d_addr_rom[  198] = 'h00000b2c; 	    wdata_rom[  198] = 'h08a5d73e; 	    wvalid_rom[  198] = 1; 
    i_addr_rom[  199] = 'h0000003c; 	    d_addr_rom[  199] = 'h00000840; 	    wdata_rom[  199] = 'h69edb675; 	    wvalid_rom[  199] = 0; 
    i_addr_rom[  200] = 'h000004d4; 	    d_addr_rom[  200] = 'h000008f4; 	    wdata_rom[  200] = 'h2684430c; 	    wvalid_rom[  200] = 0; 
    i_addr_rom[  201] = 'h00000030; 	    d_addr_rom[  201] = 'h00000910; 	    wdata_rom[  201] = 'h4bd7bea7; 	    wvalid_rom[  201] = 1; 
    i_addr_rom[  202] = 'h00000574; 	    d_addr_rom[  202] = 'h00000e58; 	    wdata_rom[  202] = 'he6f70a7b; 	    wvalid_rom[  202] = 0; 
    i_addr_rom[  203] = 'h000005f0; 	    d_addr_rom[  203] = 'h000008bc; 	    wdata_rom[  203] = 'h92922b06; 	    wvalid_rom[  203] = 1; 
    i_addr_rom[  204] = 'h00000328; 	    d_addr_rom[  204] = 'h00000c60; 	    wdata_rom[  204] = 'he968aefd; 	    wvalid_rom[  204] = 0; 
    i_addr_rom[  205] = 'h0000041c; 	    d_addr_rom[  205] = 'h00000fdc; 	    wdata_rom[  205] = 'hc51f1947; 	    wvalid_rom[  205] = 0; 
    i_addr_rom[  206] = 'h00000310; 	    d_addr_rom[  206] = 'h00000c98; 	    wdata_rom[  206] = 'hde1d0a86; 	    wvalid_rom[  206] = 1; 
    i_addr_rom[  207] = 'h000006c8; 	    d_addr_rom[  207] = 'h00000f00; 	    wdata_rom[  207] = 'h50e3c019; 	    wvalid_rom[  207] = 0; 
    i_addr_rom[  208] = 'h00000764; 	    d_addr_rom[  208] = 'h00000954; 	    wdata_rom[  208] = 'hf88e61e5; 	    wvalid_rom[  208] = 1; 
    i_addr_rom[  209] = 'h00000148; 	    d_addr_rom[  209] = 'h00000a94; 	    wdata_rom[  209] = 'hb5e33426; 	    wvalid_rom[  209] = 1; 
    i_addr_rom[  210] = 'h00000148; 	    d_addr_rom[  210] = 'h00000914; 	    wdata_rom[  210] = 'hce5aa367; 	    wvalid_rom[  210] = 1; 
    i_addr_rom[  211] = 'h00000774; 	    d_addr_rom[  211] = 'h000008b0; 	    wdata_rom[  211] = 'hae9b9058; 	    wvalid_rom[  211] = 1; 
    i_addr_rom[  212] = 'h000003b0; 	    d_addr_rom[  212] = 'h00000a20; 	    wdata_rom[  212] = 'h397dd768; 	    wvalid_rom[  212] = 1; 
    i_addr_rom[  213] = 'h00000700; 	    d_addr_rom[  213] = 'h00000bec; 	    wdata_rom[  213] = 'hea8bb25d; 	    wvalid_rom[  213] = 1; 
    i_addr_rom[  214] = 'h00000708; 	    d_addr_rom[  214] = 'h00000f68; 	    wdata_rom[  214] = 'h9dba48c0; 	    wvalid_rom[  214] = 0; 
    i_addr_rom[  215] = 'h00000528; 	    d_addr_rom[  215] = 'h00000f84; 	    wdata_rom[  215] = 'hdaac9182; 	    wvalid_rom[  215] = 1; 
    i_addr_rom[  216] = 'h00000430; 	    d_addr_rom[  216] = 'h00000c2c; 	    wdata_rom[  216] = 'h3618dbe4; 	    wvalid_rom[  216] = 0; 
    i_addr_rom[  217] = 'h000000c4; 	    d_addr_rom[  217] = 'h00000ca0; 	    wdata_rom[  217] = 'hf1aebe50; 	    wvalid_rom[  217] = 1; 
    i_addr_rom[  218] = 'h000000d4; 	    d_addr_rom[  218] = 'h00000934; 	    wdata_rom[  218] = 'h509eaace; 	    wvalid_rom[  218] = 0; 
    i_addr_rom[  219] = 'h000006c0; 	    d_addr_rom[  219] = 'h00000900; 	    wdata_rom[  219] = 'he7e6b840; 	    wvalid_rom[  219] = 1; 
    i_addr_rom[  220] = 'h0000019c; 	    d_addr_rom[  220] = 'h00000a04; 	    wdata_rom[  220] = 'h956d34c6; 	    wvalid_rom[  220] = 1; 
    i_addr_rom[  221] = 'h00000240; 	    d_addr_rom[  221] = 'h00000b48; 	    wdata_rom[  221] = 'hd8f09f1a; 	    wvalid_rom[  221] = 0; 
    i_addr_rom[  222] = 'h0000070c; 	    d_addr_rom[  222] = 'h00000f04; 	    wdata_rom[  222] = 'hc412ea85; 	    wvalid_rom[  222] = 1; 
    i_addr_rom[  223] = 'h000006c4; 	    d_addr_rom[  223] = 'h00000d44; 	    wdata_rom[  223] = 'h9907ac51; 	    wvalid_rom[  223] = 1; 
    i_addr_rom[  224] = 'h0000063c; 	    d_addr_rom[  224] = 'h00000e60; 	    wdata_rom[  224] = 'h4fbbb07e; 	    wvalid_rom[  224] = 1; 
    i_addr_rom[  225] = 'h00000158; 	    d_addr_rom[  225] = 'h0000092c; 	    wdata_rom[  225] = 'he2d20030; 	    wvalid_rom[  225] = 0; 
    i_addr_rom[  226] = 'h0000054c; 	    d_addr_rom[  226] = 'h0000080c; 	    wdata_rom[  226] = 'h227c440f; 	    wvalid_rom[  226] = 1; 
    i_addr_rom[  227] = 'h000002fc; 	    d_addr_rom[  227] = 'h00000f7c; 	    wdata_rom[  227] = 'h90ea958c; 	    wvalid_rom[  227] = 0; 
    i_addr_rom[  228] = 'h000007bc; 	    d_addr_rom[  228] = 'h00000af0; 	    wdata_rom[  228] = 'h1da0d57c; 	    wvalid_rom[  228] = 1; 
    i_addr_rom[  229] = 'h0000078c; 	    d_addr_rom[  229] = 'h00000814; 	    wdata_rom[  229] = 'h4bfc6b7f; 	    wvalid_rom[  229] = 1; 
    i_addr_rom[  230] = 'h000002b4; 	    d_addr_rom[  230] = 'h00000be8; 	    wdata_rom[  230] = 'h670b27ba; 	    wvalid_rom[  230] = 1; 
    i_addr_rom[  231] = 'h00000770; 	    d_addr_rom[  231] = 'h00000a44; 	    wdata_rom[  231] = 'h98bd2c95; 	    wvalid_rom[  231] = 0; 
    i_addr_rom[  232] = 'h000007ec; 	    d_addr_rom[  232] = 'h00000918; 	    wdata_rom[  232] = 'h7aba4bb0; 	    wvalid_rom[  232] = 0; 
    i_addr_rom[  233] = 'h000002c0; 	    d_addr_rom[  233] = 'h00000ca4; 	    wdata_rom[  233] = 'he2f70fe5; 	    wvalid_rom[  233] = 0; 
    i_addr_rom[  234] = 'h00000678; 	    d_addr_rom[  234] = 'h00000afc; 	    wdata_rom[  234] = 'h6d6e2be7; 	    wvalid_rom[  234] = 1; 
    i_addr_rom[  235] = 'h000003f0; 	    d_addr_rom[  235] = 'h00000d84; 	    wdata_rom[  235] = 'h29d9a3d5; 	    wvalid_rom[  235] = 0; 
    i_addr_rom[  236] = 'h00000494; 	    d_addr_rom[  236] = 'h00000c94; 	    wdata_rom[  236] = 'ha8637cda; 	    wvalid_rom[  236] = 1; 
    i_addr_rom[  237] = 'h0000016c; 	    d_addr_rom[  237] = 'h00000940; 	    wdata_rom[  237] = 'hab998417; 	    wvalid_rom[  237] = 1; 
    i_addr_rom[  238] = 'h0000013c; 	    d_addr_rom[  238] = 'h00000a74; 	    wdata_rom[  238] = 'h216d71a5; 	    wvalid_rom[  238] = 0; 
    i_addr_rom[  239] = 'h000004a0; 	    d_addr_rom[  239] = 'h00000ab8; 	    wdata_rom[  239] = 'hdf4ebf33; 	    wvalid_rom[  239] = 1; 
    i_addr_rom[  240] = 'h000006dc; 	    d_addr_rom[  240] = 'h00000be8; 	    wdata_rom[  240] = 'h86c008a3; 	    wvalid_rom[  240] = 1; 
    i_addr_rom[  241] = 'h000001c4; 	    d_addr_rom[  241] = 'h00000894; 	    wdata_rom[  241] = 'h9259c71a; 	    wvalid_rom[  241] = 1; 
    i_addr_rom[  242] = 'h0000079c; 	    d_addr_rom[  242] = 'h0000088c; 	    wdata_rom[  242] = 'h19641659; 	    wvalid_rom[  242] = 0; 
    i_addr_rom[  243] = 'h00000418; 	    d_addr_rom[  243] = 'h000009d4; 	    wdata_rom[  243] = 'hf8023edf; 	    wvalid_rom[  243] = 1; 
    i_addr_rom[  244] = 'h00000284; 	    d_addr_rom[  244] = 'h00000de0; 	    wdata_rom[  244] = 'h87623d90; 	    wvalid_rom[  244] = 1; 
    i_addr_rom[  245] = 'h00000440; 	    d_addr_rom[  245] = 'h00000ee0; 	    wdata_rom[  245] = 'he3f5d26d; 	    wvalid_rom[  245] = 0; 
    i_addr_rom[  246] = 'h000003a4; 	    d_addr_rom[  246] = 'h00000dec; 	    wdata_rom[  246] = 'ha445f129; 	    wvalid_rom[  246] = 1; 
    i_addr_rom[  247] = 'h00000328; 	    d_addr_rom[  247] = 'h00000850; 	    wdata_rom[  247] = 'h95af1af1; 	    wvalid_rom[  247] = 0; 
    i_addr_rom[  248] = 'h000003f0; 	    d_addr_rom[  248] = 'h00000974; 	    wdata_rom[  248] = 'hdeaa2465; 	    wvalid_rom[  248] = 1; 
    i_addr_rom[  249] = 'h00000458; 	    d_addr_rom[  249] = 'h00000d30; 	    wdata_rom[  249] = 'hb57eafc7; 	    wvalid_rom[  249] = 0; 
    i_addr_rom[  250] = 'h00000074; 	    d_addr_rom[  250] = 'h00000e98; 	    wdata_rom[  250] = 'hc6df7c34; 	    wvalid_rom[  250] = 0; 
    i_addr_rom[  251] = 'h000005d0; 	    d_addr_rom[  251] = 'h00000ed0; 	    wdata_rom[  251] = 'h6dc81922; 	    wvalid_rom[  251] = 1; 
    i_addr_rom[  252] = 'h000001c4; 	    d_addr_rom[  252] = 'h00000fa8; 	    wdata_rom[  252] = 'h0cf20fe7; 	    wvalid_rom[  252] = 1; 
    i_addr_rom[  253] = 'h000003dc; 	    d_addr_rom[  253] = 'h00000a50; 	    wdata_rom[  253] = 'hc49b63e2; 	    wvalid_rom[  253] = 1; 
    i_addr_rom[  254] = 'h000006cc; 	    d_addr_rom[  254] = 'h00000b98; 	    wdata_rom[  254] = 'h1d471687; 	    wvalid_rom[  254] = 1; 
    i_addr_rom[  255] = 'h00000100; 	    d_addr_rom[  255] = 'h00000a38; 	    wdata_rom[  255] = 'h47cc25b6; 	    wvalid_rom[  255] = 1; 
    i_addr_rom[  256] = 'h00000168; 	    d_addr_rom[  256] = 'h00000da4; 	    wdata_rom[  256] = 'he04400e5; 	    wvalid_rom[  256] = 1; 
    i_addr_rom[  257] = 'h00000080; 	    d_addr_rom[  257] = 'h00000bf8; 	    wdata_rom[  257] = 'h7b2b08fa; 	    wvalid_rom[  257] = 0; 
    i_addr_rom[  258] = 'h0000045c; 	    d_addr_rom[  258] = 'h000009c4; 	    wdata_rom[  258] = 'h5269a8af; 	    wvalid_rom[  258] = 0; 
    i_addr_rom[  259] = 'h000006d4; 	    d_addr_rom[  259] = 'h000008b8; 	    wdata_rom[  259] = 'h3d957152; 	    wvalid_rom[  259] = 1; 
    i_addr_rom[  260] = 'h00000064; 	    d_addr_rom[  260] = 'h000009a0; 	    wdata_rom[  260] = 'h9e42567b; 	    wvalid_rom[  260] = 0; 
    i_addr_rom[  261] = 'h000002c0; 	    d_addr_rom[  261] = 'h00000d6c; 	    wdata_rom[  261] = 'h39fa5897; 	    wvalid_rom[  261] = 1; 
    i_addr_rom[  262] = 'h0000026c; 	    d_addr_rom[  262] = 'h00000f7c; 	    wdata_rom[  262] = 'h0dd7753f; 	    wvalid_rom[  262] = 1; 
    i_addr_rom[  263] = 'h00000464; 	    d_addr_rom[  263] = 'h00000930; 	    wdata_rom[  263] = 'hc9937f25; 	    wvalid_rom[  263] = 1; 
    i_addr_rom[  264] = 'h00000674; 	    d_addr_rom[  264] = 'h00000fa0; 	    wdata_rom[  264] = 'hd21a7d40; 	    wvalid_rom[  264] = 1; 
    i_addr_rom[  265] = 'h00000764; 	    d_addr_rom[  265] = 'h00000fc8; 	    wdata_rom[  265] = 'h9375c834; 	    wvalid_rom[  265] = 1; 
    i_addr_rom[  266] = 'h0000016c; 	    d_addr_rom[  266] = 'h000008c0; 	    wdata_rom[  266] = 'h5c279513; 	    wvalid_rom[  266] = 1; 
    i_addr_rom[  267] = 'h0000070c; 	    d_addr_rom[  267] = 'h000009c8; 	    wdata_rom[  267] = 'hfd187170; 	    wvalid_rom[  267] = 0; 
    i_addr_rom[  268] = 'h00000144; 	    d_addr_rom[  268] = 'h00000f34; 	    wdata_rom[  268] = 'hcb2ff90a; 	    wvalid_rom[  268] = 0; 
    i_addr_rom[  269] = 'h00000040; 	    d_addr_rom[  269] = 'h00000b30; 	    wdata_rom[  269] = 'hcf3bd819; 	    wvalid_rom[  269] = 0; 
    i_addr_rom[  270] = 'h0000059c; 	    d_addr_rom[  270] = 'h000008a4; 	    wdata_rom[  270] = 'h944387ba; 	    wvalid_rom[  270] = 0; 
    i_addr_rom[  271] = 'h00000474; 	    d_addr_rom[  271] = 'h00000c7c; 	    wdata_rom[  271] = 'hf6b799c0; 	    wvalid_rom[  271] = 0; 
    i_addr_rom[  272] = 'h000004e4; 	    d_addr_rom[  272] = 'h00000c00; 	    wdata_rom[  272] = 'h50b5693b; 	    wvalid_rom[  272] = 0; 
    i_addr_rom[  273] = 'h00000130; 	    d_addr_rom[  273] = 'h00000d54; 	    wdata_rom[  273] = 'hd5f12f85; 	    wvalid_rom[  273] = 1; 
    i_addr_rom[  274] = 'h00000644; 	    d_addr_rom[  274] = 'h00000aa0; 	    wdata_rom[  274] = 'h633ef86b; 	    wvalid_rom[  274] = 0; 
    i_addr_rom[  275] = 'h00000738; 	    d_addr_rom[  275] = 'h00000be0; 	    wdata_rom[  275] = 'h1b1eb521; 	    wvalid_rom[  275] = 1; 
    i_addr_rom[  276] = 'h0000001c; 	    d_addr_rom[  276] = 'h00000828; 	    wdata_rom[  276] = 'h6db889c1; 	    wvalid_rom[  276] = 0; 
    i_addr_rom[  277] = 'h00000638; 	    d_addr_rom[  277] = 'h00000800; 	    wdata_rom[  277] = 'h892a84fa; 	    wvalid_rom[  277] = 1; 
    i_addr_rom[  278] = 'h00000238; 	    d_addr_rom[  278] = 'h00000e14; 	    wdata_rom[  278] = 'h1cf3d077; 	    wvalid_rom[  278] = 1; 
    i_addr_rom[  279] = 'h0000066c; 	    d_addr_rom[  279] = 'h00000e40; 	    wdata_rom[  279] = 'h271f218c; 	    wvalid_rom[  279] = 0; 
    i_addr_rom[  280] = 'h00000688; 	    d_addr_rom[  280] = 'h00000800; 	    wdata_rom[  280] = 'h614067f3; 	    wvalid_rom[  280] = 0; 
    i_addr_rom[  281] = 'h000002ac; 	    d_addr_rom[  281] = 'h00000e54; 	    wdata_rom[  281] = 'he14f4379; 	    wvalid_rom[  281] = 1; 
    i_addr_rom[  282] = 'h0000031c; 	    d_addr_rom[  282] = 'h00000e80; 	    wdata_rom[  282] = 'h5fc21145; 	    wvalid_rom[  282] = 0; 
    i_addr_rom[  283] = 'h0000064c; 	    d_addr_rom[  283] = 'h00000b88; 	    wdata_rom[  283] = 'hde71487e; 	    wvalid_rom[  283] = 0; 
    i_addr_rom[  284] = 'h00000134; 	    d_addr_rom[  284] = 'h00000d60; 	    wdata_rom[  284] = 'h9a941f69; 	    wvalid_rom[  284] = 1; 
    i_addr_rom[  285] = 'h00000538; 	    d_addr_rom[  285] = 'h00000d58; 	    wdata_rom[  285] = 'h2c954295; 	    wvalid_rom[  285] = 0; 
    i_addr_rom[  286] = 'h00000530; 	    d_addr_rom[  286] = 'h00000984; 	    wdata_rom[  286] = 'he9f08043; 	    wvalid_rom[  286] = 1; 
    i_addr_rom[  287] = 'h00000734; 	    d_addr_rom[  287] = 'h00000b54; 	    wdata_rom[  287] = 'hf0e56080; 	    wvalid_rom[  287] = 0; 
    i_addr_rom[  288] = 'h000000bc; 	    d_addr_rom[  288] = 'h000008e0; 	    wdata_rom[  288] = 'hc4eaaa48; 	    wvalid_rom[  288] = 1; 
    i_addr_rom[  289] = 'h00000474; 	    d_addr_rom[  289] = 'h00000e20; 	    wdata_rom[  289] = 'h26bdd1a0; 	    wvalid_rom[  289] = 0; 
    i_addr_rom[  290] = 'h00000158; 	    d_addr_rom[  290] = 'h00000fb8; 	    wdata_rom[  290] = 'h924f806c; 	    wvalid_rom[  290] = 1; 
    i_addr_rom[  291] = 'h00000630; 	    d_addr_rom[  291] = 'h00000a5c; 	    wdata_rom[  291] = 'he692fbda; 	    wvalid_rom[  291] = 1; 
    i_addr_rom[  292] = 'h0000074c; 	    d_addr_rom[  292] = 'h00000bd4; 	    wdata_rom[  292] = 'hbcc21461; 	    wvalid_rom[  292] = 1; 
    i_addr_rom[  293] = 'h00000388; 	    d_addr_rom[  293] = 'h00000df4; 	    wdata_rom[  293] = 'hea891c44; 	    wvalid_rom[  293] = 0; 
    i_addr_rom[  294] = 'h000000d8; 	    d_addr_rom[  294] = 'h00000c44; 	    wdata_rom[  294] = 'h4a1afaae; 	    wvalid_rom[  294] = 0; 
    i_addr_rom[  295] = 'h00000654; 	    d_addr_rom[  295] = 'h00000cac; 	    wdata_rom[  295] = 'h71fb5479; 	    wvalid_rom[  295] = 1; 
    i_addr_rom[  296] = 'h0000049c; 	    d_addr_rom[  296] = 'h00000fb0; 	    wdata_rom[  296] = 'h05a912ae; 	    wvalid_rom[  296] = 0; 
    i_addr_rom[  297] = 'h000002f4; 	    d_addr_rom[  297] = 'h00000bac; 	    wdata_rom[  297] = 'h20749344; 	    wvalid_rom[  297] = 0; 
    i_addr_rom[  298] = 'h0000049c; 	    d_addr_rom[  298] = 'h00000aa0; 	    wdata_rom[  298] = 'h6e2c7784; 	    wvalid_rom[  298] = 0; 
    i_addr_rom[  299] = 'h000003c8; 	    d_addr_rom[  299] = 'h00000b24; 	    wdata_rom[  299] = 'h11f01f38; 	    wvalid_rom[  299] = 0; 
    i_addr_rom[  300] = 'h000001dc; 	    d_addr_rom[  300] = 'h00000cd0; 	    wdata_rom[  300] = 'h9c6c78cf; 	    wvalid_rom[  300] = 1; 
    i_addr_rom[  301] = 'h00000348; 	    d_addr_rom[  301] = 'h00000ca4; 	    wdata_rom[  301] = 'hc1f4e19d; 	    wvalid_rom[  301] = 0; 
    i_addr_rom[  302] = 'h0000008c; 	    d_addr_rom[  302] = 'h00000af0; 	    wdata_rom[  302] = 'hdc885977; 	    wvalid_rom[  302] = 1; 
    i_addr_rom[  303] = 'h000003e8; 	    d_addr_rom[  303] = 'h00000c58; 	    wdata_rom[  303] = 'h0fd1d46e; 	    wvalid_rom[  303] = 1; 
    i_addr_rom[  304] = 'h0000057c; 	    d_addr_rom[  304] = 'h000008d4; 	    wdata_rom[  304] = 'h88afba5c; 	    wvalid_rom[  304] = 1; 
    i_addr_rom[  305] = 'h00000288; 	    d_addr_rom[  305] = 'h00000958; 	    wdata_rom[  305] = 'h19c8706d; 	    wvalid_rom[  305] = 1; 
    i_addr_rom[  306] = 'h0000050c; 	    d_addr_rom[  306] = 'h00000ee0; 	    wdata_rom[  306] = 'h8912c4cd; 	    wvalid_rom[  306] = 1; 
    i_addr_rom[  307] = 'h00000674; 	    d_addr_rom[  307] = 'h00000fc0; 	    wdata_rom[  307] = 'h363e773d; 	    wvalid_rom[  307] = 1; 
    i_addr_rom[  308] = 'h00000644; 	    d_addr_rom[  308] = 'h00000c60; 	    wdata_rom[  308] = 'h13958272; 	    wvalid_rom[  308] = 0; 
    i_addr_rom[  309] = 'h00000604; 	    d_addr_rom[  309] = 'h00000f70; 	    wdata_rom[  309] = 'h1845b7e1; 	    wvalid_rom[  309] = 1; 
    i_addr_rom[  310] = 'h000000d4; 	    d_addr_rom[  310] = 'h00000d70; 	    wdata_rom[  310] = 'had6b4933; 	    wvalid_rom[  310] = 0; 
    i_addr_rom[  311] = 'h0000019c; 	    d_addr_rom[  311] = 'h000008d0; 	    wdata_rom[  311] = 'h935a3498; 	    wvalid_rom[  311] = 0; 
    i_addr_rom[  312] = 'h000004ac; 	    d_addr_rom[  312] = 'h00000af8; 	    wdata_rom[  312] = 'h45bcca37; 	    wvalid_rom[  312] = 0; 
    i_addr_rom[  313] = 'h00000384; 	    d_addr_rom[  313] = 'h00000bc8; 	    wdata_rom[  313] = 'h2332240e; 	    wvalid_rom[  313] = 0; 
    i_addr_rom[  314] = 'h00000398; 	    d_addr_rom[  314] = 'h00000e78; 	    wdata_rom[  314] = 'hc2220736; 	    wvalid_rom[  314] = 0; 
    i_addr_rom[  315] = 'h000002c8; 	    d_addr_rom[  315] = 'h00000b18; 	    wdata_rom[  315] = 'hd0c82ab3; 	    wvalid_rom[  315] = 1; 
    i_addr_rom[  316] = 'h0000006c; 	    d_addr_rom[  316] = 'h00000920; 	    wdata_rom[  316] = 'ha4bcd6dc; 	    wvalid_rom[  316] = 0; 
    i_addr_rom[  317] = 'h0000040c; 	    d_addr_rom[  317] = 'h00000f90; 	    wdata_rom[  317] = 'hb271de18; 	    wvalid_rom[  317] = 1; 
    i_addr_rom[  318] = 'h0000003c; 	    d_addr_rom[  318] = 'h00000b30; 	    wdata_rom[  318] = 'hebc623ee; 	    wvalid_rom[  318] = 0; 
    i_addr_rom[  319] = 'h00000368; 	    d_addr_rom[  319] = 'h00000c6c; 	    wdata_rom[  319] = 'hdd61c0f8; 	    wvalid_rom[  319] = 1; 
    i_addr_rom[  320] = 'h00000278; 	    d_addr_rom[  320] = 'h00000db8; 	    wdata_rom[  320] = 'h42514a64; 	    wvalid_rom[  320] = 1; 
    i_addr_rom[  321] = 'h00000724; 	    d_addr_rom[  321] = 'h0000080c; 	    wdata_rom[  321] = 'h31b86e90; 	    wvalid_rom[  321] = 0; 
    i_addr_rom[  322] = 'h000004a0; 	    d_addr_rom[  322] = 'h00000fdc; 	    wdata_rom[  322] = 'hdf386c1e; 	    wvalid_rom[  322] = 1; 
    i_addr_rom[  323] = 'h000006ec; 	    d_addr_rom[  323] = 'h00000b80; 	    wdata_rom[  323] = 'h81822bbd; 	    wvalid_rom[  323] = 0; 
    i_addr_rom[  324] = 'h00000168; 	    d_addr_rom[  324] = 'h00000be0; 	    wdata_rom[  324] = 'he64a09d8; 	    wvalid_rom[  324] = 0; 
    i_addr_rom[  325] = 'h00000654; 	    d_addr_rom[  325] = 'h00000ccc; 	    wdata_rom[  325] = 'h41716525; 	    wvalid_rom[  325] = 1; 
    i_addr_rom[  326] = 'h00000660; 	    d_addr_rom[  326] = 'h00000e38; 	    wdata_rom[  326] = 'h72b72733; 	    wvalid_rom[  326] = 0; 
    i_addr_rom[  327] = 'h00000638; 	    d_addr_rom[  327] = 'h00000af0; 	    wdata_rom[  327] = 'ha35bd143; 	    wvalid_rom[  327] = 0; 
    i_addr_rom[  328] = 'h0000070c; 	    d_addr_rom[  328] = 'h00000f3c; 	    wdata_rom[  328] = 'ha072e18b; 	    wvalid_rom[  328] = 0; 
    i_addr_rom[  329] = 'h00000410; 	    d_addr_rom[  329] = 'h00000f10; 	    wdata_rom[  329] = 'h038d44db; 	    wvalid_rom[  329] = 1; 
    i_addr_rom[  330] = 'h000002c4; 	    d_addr_rom[  330] = 'h00000c8c; 	    wdata_rom[  330] = 'hd2ee1ad4; 	    wvalid_rom[  330] = 1; 
    i_addr_rom[  331] = 'h000007a4; 	    d_addr_rom[  331] = 'h0000083c; 	    wdata_rom[  331] = 'hf3ca5ea5; 	    wvalid_rom[  331] = 1; 
    i_addr_rom[  332] = 'h00000644; 	    d_addr_rom[  332] = 'h00000bf8; 	    wdata_rom[  332] = 'h2c4121c8; 	    wvalid_rom[  332] = 1; 
    i_addr_rom[  333] = 'h0000062c; 	    d_addr_rom[  333] = 'h00000d30; 	    wdata_rom[  333] = 'h63cf7333; 	    wvalid_rom[  333] = 1; 
    i_addr_rom[  334] = 'h000005cc; 	    d_addr_rom[  334] = 'h00000f08; 	    wdata_rom[  334] = 'h2476d93e; 	    wvalid_rom[  334] = 1; 
    i_addr_rom[  335] = 'h00000438; 	    d_addr_rom[  335] = 'h00000aec; 	    wdata_rom[  335] = 'h46845232; 	    wvalid_rom[  335] = 1; 
    i_addr_rom[  336] = 'h000005b0; 	    d_addr_rom[  336] = 'h00000c1c; 	    wdata_rom[  336] = 'h13d9ca42; 	    wvalid_rom[  336] = 0; 
    i_addr_rom[  337] = 'h0000001c; 	    d_addr_rom[  337] = 'h00000868; 	    wdata_rom[  337] = 'h93ab566a; 	    wvalid_rom[  337] = 1; 
    i_addr_rom[  338] = 'h00000444; 	    d_addr_rom[  338] = 'h00000d20; 	    wdata_rom[  338] = 'h1fad7327; 	    wvalid_rom[  338] = 0; 
    i_addr_rom[  339] = 'h000003a8; 	    d_addr_rom[  339] = 'h00000d78; 	    wdata_rom[  339] = 'h1ef544c8; 	    wvalid_rom[  339] = 1; 
    i_addr_rom[  340] = 'h0000027c; 	    d_addr_rom[  340] = 'h00000fa0; 	    wdata_rom[  340] = 'h9df924f0; 	    wvalid_rom[  340] = 1; 
    i_addr_rom[  341] = 'h000002e0; 	    d_addr_rom[  341] = 'h000008c4; 	    wdata_rom[  341] = 'h0332499f; 	    wvalid_rom[  341] = 0; 
    i_addr_rom[  342] = 'h00000348; 	    d_addr_rom[  342] = 'h00000e04; 	    wdata_rom[  342] = 'h14cee293; 	    wvalid_rom[  342] = 1; 
    i_addr_rom[  343] = 'h00000234; 	    d_addr_rom[  343] = 'h00000a84; 	    wdata_rom[  343] = 'hd104e2bc; 	    wvalid_rom[  343] = 0; 
    i_addr_rom[  344] = 'h000002f0; 	    d_addr_rom[  344] = 'h00000ee8; 	    wdata_rom[  344] = 'h7d274047; 	    wvalid_rom[  344] = 1; 
    i_addr_rom[  345] = 'h000006d8; 	    d_addr_rom[  345] = 'h00000b0c; 	    wdata_rom[  345] = 'h47d0b412; 	    wvalid_rom[  345] = 0; 
    i_addr_rom[  346] = 'h00000210; 	    d_addr_rom[  346] = 'h00000d10; 	    wdata_rom[  346] = 'ha94c73f9; 	    wvalid_rom[  346] = 0; 
    i_addr_rom[  347] = 'h000005ac; 	    d_addr_rom[  347] = 'h00000ef8; 	    wdata_rom[  347] = 'h9048324b; 	    wvalid_rom[  347] = 0; 
    i_addr_rom[  348] = 'h0000046c; 	    d_addr_rom[  348] = 'h00000a20; 	    wdata_rom[  348] = 'h81d06ba8; 	    wvalid_rom[  348] = 0; 
    i_addr_rom[  349] = 'h000007c4; 	    d_addr_rom[  349] = 'h00000c78; 	    wdata_rom[  349] = 'he2380053; 	    wvalid_rom[  349] = 1; 
    i_addr_rom[  350] = 'h00000088; 	    d_addr_rom[  350] = 'h00000d74; 	    wdata_rom[  350] = 'h5f385f90; 	    wvalid_rom[  350] = 0; 
    i_addr_rom[  351] = 'h000007e0; 	    d_addr_rom[  351] = 'h00000a04; 	    wdata_rom[  351] = 'h1a7d9a5b; 	    wvalid_rom[  351] = 0; 
    i_addr_rom[  352] = 'h00000310; 	    d_addr_rom[  352] = 'h00000ff8; 	    wdata_rom[  352] = 'h8c95beac; 	    wvalid_rom[  352] = 1; 
    i_addr_rom[  353] = 'h000003f8; 	    d_addr_rom[  353] = 'h00000d48; 	    wdata_rom[  353] = 'h1c5e5bed; 	    wvalid_rom[  353] = 1; 
    i_addr_rom[  354] = 'h00000328; 	    d_addr_rom[  354] = 'h000009ec; 	    wdata_rom[  354] = 'h1f3b7bfa; 	    wvalid_rom[  354] = 1; 
    i_addr_rom[  355] = 'h000000a4; 	    d_addr_rom[  355] = 'h00000fe8; 	    wdata_rom[  355] = 'h93b981b2; 	    wvalid_rom[  355] = 0; 
    i_addr_rom[  356] = 'h000007cc; 	    d_addr_rom[  356] = 'h00000ec4; 	    wdata_rom[  356] = 'h17eeefa7; 	    wvalid_rom[  356] = 0; 
    i_addr_rom[  357] = 'h00000738; 	    d_addr_rom[  357] = 'h00000f48; 	    wdata_rom[  357] = 'h1fb22e06; 	    wvalid_rom[  357] = 0; 
    i_addr_rom[  358] = 'h000000f4; 	    d_addr_rom[  358] = 'h00000940; 	    wdata_rom[  358] = 'h795b88f4; 	    wvalid_rom[  358] = 1; 
    i_addr_rom[  359] = 'h000000dc; 	    d_addr_rom[  359] = 'h000009b8; 	    wdata_rom[  359] = 'h518da9b0; 	    wvalid_rom[  359] = 1; 
    i_addr_rom[  360] = 'h00000178; 	    d_addr_rom[  360] = 'h00000eec; 	    wdata_rom[  360] = 'he955bfef; 	    wvalid_rom[  360] = 1; 
    i_addr_rom[  361] = 'h00000634; 	    d_addr_rom[  361] = 'h00000e84; 	    wdata_rom[  361] = 'hd76e2d17; 	    wvalid_rom[  361] = 1; 
    i_addr_rom[  362] = 'h0000066c; 	    d_addr_rom[  362] = 'h00000acc; 	    wdata_rom[  362] = 'hc9b0d8be; 	    wvalid_rom[  362] = 0; 
    i_addr_rom[  363] = 'h00000028; 	    d_addr_rom[  363] = 'h00000f60; 	    wdata_rom[  363] = 'hd874d169; 	    wvalid_rom[  363] = 1; 
    i_addr_rom[  364] = 'h00000254; 	    d_addr_rom[  364] = 'h000009f8; 	    wdata_rom[  364] = 'h36f9ec78; 	    wvalid_rom[  364] = 1; 
    i_addr_rom[  365] = 'h000003a8; 	    d_addr_rom[  365] = 'h00000840; 	    wdata_rom[  365] = 'h69708aee; 	    wvalid_rom[  365] = 1; 
    i_addr_rom[  366] = 'h000000b0; 	    d_addr_rom[  366] = 'h00000f3c; 	    wdata_rom[  366] = 'h022b169d; 	    wvalid_rom[  366] = 1; 
    i_addr_rom[  367] = 'h00000708; 	    d_addr_rom[  367] = 'h00000d54; 	    wdata_rom[  367] = 'h8e6ec3e7; 	    wvalid_rom[  367] = 0; 
    i_addr_rom[  368] = 'h000005a4; 	    d_addr_rom[  368] = 'h000009a4; 	    wdata_rom[  368] = 'hd8483ab1; 	    wvalid_rom[  368] = 1; 
    i_addr_rom[  369] = 'h00000510; 	    d_addr_rom[  369] = 'h00000c90; 	    wdata_rom[  369] = 'ha8649215; 	    wvalid_rom[  369] = 0; 
    i_addr_rom[  370] = 'h000007d8; 	    d_addr_rom[  370] = 'h00000b58; 	    wdata_rom[  370] = 'he11b746a; 	    wvalid_rom[  370] = 1; 
    i_addr_rom[  371] = 'h000006f4; 	    d_addr_rom[  371] = 'h00000c74; 	    wdata_rom[  371] = 'h0a1a5a84; 	    wvalid_rom[  371] = 1; 
    i_addr_rom[  372] = 'h00000740; 	    d_addr_rom[  372] = 'h00000944; 	    wdata_rom[  372] = 'h7d8ca585; 	    wvalid_rom[  372] = 1; 
    i_addr_rom[  373] = 'h00000080; 	    d_addr_rom[  373] = 'h00000bec; 	    wdata_rom[  373] = 'hbc86c428; 	    wvalid_rom[  373] = 1; 
    i_addr_rom[  374] = 'h00000340; 	    d_addr_rom[  374] = 'h00000d50; 	    wdata_rom[  374] = 'hc348a944; 	    wvalid_rom[  374] = 0; 
    i_addr_rom[  375] = 'h000006bc; 	    d_addr_rom[  375] = 'h00000c38; 	    wdata_rom[  375] = 'h521aa55d; 	    wvalid_rom[  375] = 1; 
    i_addr_rom[  376] = 'h00000538; 	    d_addr_rom[  376] = 'h0000094c; 	    wdata_rom[  376] = 'h5acec3f9; 	    wvalid_rom[  376] = 1; 
    i_addr_rom[  377] = 'h000000cc; 	    d_addr_rom[  377] = 'h00000910; 	    wdata_rom[  377] = 'hf5e9cfe6; 	    wvalid_rom[  377] = 1; 
    i_addr_rom[  378] = 'h00000150; 	    d_addr_rom[  378] = 'h00000fcc; 	    wdata_rom[  378] = 'hf0627232; 	    wvalid_rom[  378] = 1; 
    i_addr_rom[  379] = 'h00000168; 	    d_addr_rom[  379] = 'h00000c38; 	    wdata_rom[  379] = 'hc5112923; 	    wvalid_rom[  379] = 1; 
    i_addr_rom[  380] = 'h000002f0; 	    d_addr_rom[  380] = 'h00000d68; 	    wdata_rom[  380] = 'h36c70252; 	    wvalid_rom[  380] = 1; 
    i_addr_rom[  381] = 'h00000738; 	    d_addr_rom[  381] = 'h00000f70; 	    wdata_rom[  381] = 'h7e297fca; 	    wvalid_rom[  381] = 1; 
    i_addr_rom[  382] = 'h000001dc; 	    d_addr_rom[  382] = 'h00000a00; 	    wdata_rom[  382] = 'h8c8ddd77; 	    wvalid_rom[  382] = 1; 
    i_addr_rom[  383] = 'h000000f4; 	    d_addr_rom[  383] = 'h00000e50; 	    wdata_rom[  383] = 'h36ac496e; 	    wvalid_rom[  383] = 0; 
    i_addr_rom[  384] = 'h00000168; 	    d_addr_rom[  384] = 'h00000f88; 	    wdata_rom[  384] = 'h27270ad3; 	    wvalid_rom[  384] = 1; 
    i_addr_rom[  385] = 'h00000770; 	    d_addr_rom[  385] = 'h00000c60; 	    wdata_rom[  385] = 'h180ad4dd; 	    wvalid_rom[  385] = 0; 
    i_addr_rom[  386] = 'h0000076c; 	    d_addr_rom[  386] = 'h00000ce8; 	    wdata_rom[  386] = 'h44c9fe25; 	    wvalid_rom[  386] = 0; 
    i_addr_rom[  387] = 'h000003a8; 	    d_addr_rom[  387] = 'h000008f0; 	    wdata_rom[  387] = 'h736bc6ad; 	    wvalid_rom[  387] = 1; 
    i_addr_rom[  388] = 'h00000078; 	    d_addr_rom[  388] = 'h00000bf0; 	    wdata_rom[  388] = 'h9b091465; 	    wvalid_rom[  388] = 0; 
    i_addr_rom[  389] = 'h00000700; 	    d_addr_rom[  389] = 'h00000bec; 	    wdata_rom[  389] = 'h1792372a; 	    wvalid_rom[  389] = 1; 
    i_addr_rom[  390] = 'h000007b4; 	    d_addr_rom[  390] = 'h00000f1c; 	    wdata_rom[  390] = 'hd491e68c; 	    wvalid_rom[  390] = 0; 
    i_addr_rom[  391] = 'h00000194; 	    d_addr_rom[  391] = 'h00000868; 	    wdata_rom[  391] = 'h65788f50; 	    wvalid_rom[  391] = 1; 
    i_addr_rom[  392] = 'h00000324; 	    d_addr_rom[  392] = 'h00000b5c; 	    wdata_rom[  392] = 'h3eccd330; 	    wvalid_rom[  392] = 0; 
    i_addr_rom[  393] = 'h000007a4; 	    d_addr_rom[  393] = 'h00000d60; 	    wdata_rom[  393] = 'h08d4702a; 	    wvalid_rom[  393] = 0; 
    i_addr_rom[  394] = 'h00000748; 	    d_addr_rom[  394] = 'h00000eb8; 	    wdata_rom[  394] = 'h71ab8318; 	    wvalid_rom[  394] = 0; 
    i_addr_rom[  395] = 'h000006c0; 	    d_addr_rom[  395] = 'h0000088c; 	    wdata_rom[  395] = 'hd043e50f; 	    wvalid_rom[  395] = 1; 
    i_addr_rom[  396] = 'h0000024c; 	    d_addr_rom[  396] = 'h00000b98; 	    wdata_rom[  396] = 'h1a6c7b83; 	    wvalid_rom[  396] = 0; 
    i_addr_rom[  397] = 'h000001e0; 	    d_addr_rom[  397] = 'h00000da0; 	    wdata_rom[  397] = 'h3028ed89; 	    wvalid_rom[  397] = 0; 
    i_addr_rom[  398] = 'h000006f8; 	    d_addr_rom[  398] = 'h00000dc8; 	    wdata_rom[  398] = 'h651bfe6c; 	    wvalid_rom[  398] = 0; 
    i_addr_rom[  399] = 'h00000294; 	    d_addr_rom[  399] = 'h00000eb0; 	    wdata_rom[  399] = 'hc25906ee; 	    wvalid_rom[  399] = 1; 
    i_addr_rom[  400] = 'h000000d8; 	    d_addr_rom[  400] = 'h00000d18; 	    wdata_rom[  400] = 'h2f735b8f; 	    wvalid_rom[  400] = 1; 
    i_addr_rom[  401] = 'h000002c0; 	    d_addr_rom[  401] = 'h000008f4; 	    wdata_rom[  401] = 'h2c9f4e77; 	    wvalid_rom[  401] = 0; 
    i_addr_rom[  402] = 'h0000005c; 	    d_addr_rom[  402] = 'h00000fc8; 	    wdata_rom[  402] = 'hcf55d53a; 	    wvalid_rom[  402] = 0; 
    i_addr_rom[  403] = 'h00000344; 	    d_addr_rom[  403] = 'h00000844; 	    wdata_rom[  403] = 'h3fc0f39e; 	    wvalid_rom[  403] = 0; 
    i_addr_rom[  404] = 'h000003ec; 	    d_addr_rom[  404] = 'h00000d74; 	    wdata_rom[  404] = 'hdb599239; 	    wvalid_rom[  404] = 0; 
    i_addr_rom[  405] = 'h000007d8; 	    d_addr_rom[  405] = 'h00000888; 	    wdata_rom[  405] = 'hdb2c9bbe; 	    wvalid_rom[  405] = 0; 
    i_addr_rom[  406] = 'h0000017c; 	    d_addr_rom[  406] = 'h0000099c; 	    wdata_rom[  406] = 'h0d395539; 	    wvalid_rom[  406] = 0; 
    i_addr_rom[  407] = 'h00000498; 	    d_addr_rom[  407] = 'h00000e40; 	    wdata_rom[  407] = 'h7bd2df10; 	    wvalid_rom[  407] = 1; 
    i_addr_rom[  408] = 'h000005b0; 	    d_addr_rom[  408] = 'h0000099c; 	    wdata_rom[  408] = 'h8b249d25; 	    wvalid_rom[  408] = 0; 
    i_addr_rom[  409] = 'h00000564; 	    d_addr_rom[  409] = 'h00000880; 	    wdata_rom[  409] = 'h46e3375d; 	    wvalid_rom[  409] = 0; 
    i_addr_rom[  410] = 'h000005a8; 	    d_addr_rom[  410] = 'h00000dc8; 	    wdata_rom[  410] = 'haa5fc0e3; 	    wvalid_rom[  410] = 0; 
    i_addr_rom[  411] = 'h00000028; 	    d_addr_rom[  411] = 'h00000dbc; 	    wdata_rom[  411] = 'h92bc7014; 	    wvalid_rom[  411] = 0; 
    i_addr_rom[  412] = 'h00000364; 	    d_addr_rom[  412] = 'h00000d80; 	    wdata_rom[  412] = 'h007bdab5; 	    wvalid_rom[  412] = 0; 
    i_addr_rom[  413] = 'h000007c8; 	    d_addr_rom[  413] = 'h0000089c; 	    wdata_rom[  413] = 'hdae15dcc; 	    wvalid_rom[  413] = 0; 
    i_addr_rom[  414] = 'h00000144; 	    d_addr_rom[  414] = 'h00000e40; 	    wdata_rom[  414] = 'hb8629fbb; 	    wvalid_rom[  414] = 1; 
    i_addr_rom[  415] = 'h0000024c; 	    d_addr_rom[  415] = 'h000009fc; 	    wdata_rom[  415] = 'h73ceffb2; 	    wvalid_rom[  415] = 0; 
    i_addr_rom[  416] = 'h00000104; 	    d_addr_rom[  416] = 'h000008ac; 	    wdata_rom[  416] = 'h073846e6; 	    wvalid_rom[  416] = 1; 
    i_addr_rom[  417] = 'h00000470; 	    d_addr_rom[  417] = 'h00000f8c; 	    wdata_rom[  417] = 'h4f6bca62; 	    wvalid_rom[  417] = 1; 
    i_addr_rom[  418] = 'h00000484; 	    d_addr_rom[  418] = 'h00000eb8; 	    wdata_rom[  418] = 'h026fcfa6; 	    wvalid_rom[  418] = 1; 
    i_addr_rom[  419] = 'h00000054; 	    d_addr_rom[  419] = 'h00000e98; 	    wdata_rom[  419] = 'hf86110b3; 	    wvalid_rom[  419] = 0; 
    i_addr_rom[  420] = 'h0000021c; 	    d_addr_rom[  420] = 'h00000c34; 	    wdata_rom[  420] = 'h064531be; 	    wvalid_rom[  420] = 1; 
    i_addr_rom[  421] = 'h000000c0; 	    d_addr_rom[  421] = 'h0000085c; 	    wdata_rom[  421] = 'h9cdd81b5; 	    wvalid_rom[  421] = 0; 
    i_addr_rom[  422] = 'h000005c4; 	    d_addr_rom[  422] = 'h00000d30; 	    wdata_rom[  422] = 'hcf817bb8; 	    wvalid_rom[  422] = 1; 
    i_addr_rom[  423] = 'h00000614; 	    d_addr_rom[  423] = 'h00000ae4; 	    wdata_rom[  423] = 'h27b48f4d; 	    wvalid_rom[  423] = 0; 
    i_addr_rom[  424] = 'h00000788; 	    d_addr_rom[  424] = 'h00000b24; 	    wdata_rom[  424] = 'h084e92d3; 	    wvalid_rom[  424] = 0; 
    i_addr_rom[  425] = 'h00000450; 	    d_addr_rom[  425] = 'h00000d7c; 	    wdata_rom[  425] = 'h94f54e00; 	    wvalid_rom[  425] = 1; 
    i_addr_rom[  426] = 'h00000724; 	    d_addr_rom[  426] = 'h00000e44; 	    wdata_rom[  426] = 'hecec3968; 	    wvalid_rom[  426] = 1; 
    i_addr_rom[  427] = 'h00000614; 	    d_addr_rom[  427] = 'h000009d8; 	    wdata_rom[  427] = 'hb722f593; 	    wvalid_rom[  427] = 0; 
    i_addr_rom[  428] = 'h000007a4; 	    d_addr_rom[  428] = 'h00000e84; 	    wdata_rom[  428] = 'h1fff4289; 	    wvalid_rom[  428] = 1; 
    i_addr_rom[  429] = 'h000003c8; 	    d_addr_rom[  429] = 'h00000f50; 	    wdata_rom[  429] = 'h0da32349; 	    wvalid_rom[  429] = 0; 
    i_addr_rom[  430] = 'h0000015c; 	    d_addr_rom[  430] = 'h00000e78; 	    wdata_rom[  430] = 'h6e4bbc44; 	    wvalid_rom[  430] = 0; 
    i_addr_rom[  431] = 'h000006e0; 	    d_addr_rom[  431] = 'h000008a4; 	    wdata_rom[  431] = 'hf61aeef6; 	    wvalid_rom[  431] = 0; 
    i_addr_rom[  432] = 'h000001d4; 	    d_addr_rom[  432] = 'h00000bd4; 	    wdata_rom[  432] = 'h36ad50b7; 	    wvalid_rom[  432] = 0; 
    i_addr_rom[  433] = 'h000002dc; 	    d_addr_rom[  433] = 'h00000f94; 	    wdata_rom[  433] = 'h419ceb4a; 	    wvalid_rom[  433] = 1; 
    i_addr_rom[  434] = 'h00000050; 	    d_addr_rom[  434] = 'h00000814; 	    wdata_rom[  434] = 'h0d182a29; 	    wvalid_rom[  434] = 0; 
    i_addr_rom[  435] = 'h00000228; 	    d_addr_rom[  435] = 'h00000bcc; 	    wdata_rom[  435] = 'h832a5660; 	    wvalid_rom[  435] = 1; 
    i_addr_rom[  436] = 'h00000364; 	    d_addr_rom[  436] = 'h00000d48; 	    wdata_rom[  436] = 'h957a6748; 	    wvalid_rom[  436] = 0; 
    i_addr_rom[  437] = 'h000000cc; 	    d_addr_rom[  437] = 'h000009ac; 	    wdata_rom[  437] = 'h30e77323; 	    wvalid_rom[  437] = 0; 
    i_addr_rom[  438] = 'h00000510; 	    d_addr_rom[  438] = 'h00000ac8; 	    wdata_rom[  438] = 'hb839157e; 	    wvalid_rom[  438] = 0; 
    i_addr_rom[  439] = 'h0000057c; 	    d_addr_rom[  439] = 'h00000f94; 	    wdata_rom[  439] = 'ha2dbc430; 	    wvalid_rom[  439] = 1; 
    i_addr_rom[  440] = 'h00000678; 	    d_addr_rom[  440] = 'h00000974; 	    wdata_rom[  440] = 'h4adf51e7; 	    wvalid_rom[  440] = 1; 
    i_addr_rom[  441] = 'h000000e4; 	    d_addr_rom[  441] = 'h0000096c; 	    wdata_rom[  441] = 'ha19e59f3; 	    wvalid_rom[  441] = 1; 
    i_addr_rom[  442] = 'h00000300; 	    d_addr_rom[  442] = 'h00000a50; 	    wdata_rom[  442] = 'h90f327a2; 	    wvalid_rom[  442] = 0; 
    i_addr_rom[  443] = 'h00000270; 	    d_addr_rom[  443] = 'h00000d6c; 	    wdata_rom[  443] = 'h51757757; 	    wvalid_rom[  443] = 0; 
    i_addr_rom[  444] = 'h00000080; 	    d_addr_rom[  444] = 'h00000b28; 	    wdata_rom[  444] = 'h6a041b15; 	    wvalid_rom[  444] = 0; 
    i_addr_rom[  445] = 'h000001e0; 	    d_addr_rom[  445] = 'h00000ea0; 	    wdata_rom[  445] = 'h461cd112; 	    wvalid_rom[  445] = 0; 
    i_addr_rom[  446] = 'h000007dc; 	    d_addr_rom[  446] = 'h00000e3c; 	    wdata_rom[  446] = 'hb2b654a6; 	    wvalid_rom[  446] = 1; 
    i_addr_rom[  447] = 'h00000558; 	    d_addr_rom[  447] = 'h00000fd4; 	    wdata_rom[  447] = 'h3460d19c; 	    wvalid_rom[  447] = 0; 
    i_addr_rom[  448] = 'h000000dc; 	    d_addr_rom[  448] = 'h00000b54; 	    wdata_rom[  448] = 'h20969397; 	    wvalid_rom[  448] = 0; 
    i_addr_rom[  449] = 'h0000000c; 	    d_addr_rom[  449] = 'h00000ec8; 	    wdata_rom[  449] = 'hc6c4ad73; 	    wvalid_rom[  449] = 0; 
    i_addr_rom[  450] = 'h0000017c; 	    d_addr_rom[  450] = 'h00000e94; 	    wdata_rom[  450] = 'h7ff9a550; 	    wvalid_rom[  450] = 1; 
    i_addr_rom[  451] = 'h000007bc; 	    d_addr_rom[  451] = 'h0000084c; 	    wdata_rom[  451] = 'h75cfebc4; 	    wvalid_rom[  451] = 0; 
    i_addr_rom[  452] = 'h000000fc; 	    d_addr_rom[  452] = 'h00000c3c; 	    wdata_rom[  452] = 'h37db2094; 	    wvalid_rom[  452] = 0; 
    i_addr_rom[  453] = 'h000005c8; 	    d_addr_rom[  453] = 'h00000e54; 	    wdata_rom[  453] = 'h06399952; 	    wvalid_rom[  453] = 0; 
    i_addr_rom[  454] = 'h00000730; 	    d_addr_rom[  454] = 'h00000aac; 	    wdata_rom[  454] = 'h1607ee36; 	    wvalid_rom[  454] = 1; 
    i_addr_rom[  455] = 'h0000048c; 	    d_addr_rom[  455] = 'h00000cac; 	    wdata_rom[  455] = 'he140f9a7; 	    wvalid_rom[  455] = 1; 
    i_addr_rom[  456] = 'h00000468; 	    d_addr_rom[  456] = 'h00000edc; 	    wdata_rom[  456] = 'h67146f13; 	    wvalid_rom[  456] = 1; 
    i_addr_rom[  457] = 'h000003d0; 	    d_addr_rom[  457] = 'h00000d8c; 	    wdata_rom[  457] = 'hd6b99eb3; 	    wvalid_rom[  457] = 1; 
    i_addr_rom[  458] = 'h00000458; 	    d_addr_rom[  458] = 'h00000e3c; 	    wdata_rom[  458] = 'h17eb9937; 	    wvalid_rom[  458] = 0; 
    i_addr_rom[  459] = 'h000001a8; 	    d_addr_rom[  459] = 'h00000b9c; 	    wdata_rom[  459] = 'hf110b229; 	    wvalid_rom[  459] = 0; 
    i_addr_rom[  460] = 'h000004bc; 	    d_addr_rom[  460] = 'h00000be0; 	    wdata_rom[  460] = 'h51a9a83d; 	    wvalid_rom[  460] = 0; 
    i_addr_rom[  461] = 'h000005c4; 	    d_addr_rom[  461] = 'h000009e0; 	    wdata_rom[  461] = 'he52ba4db; 	    wvalid_rom[  461] = 1; 
    i_addr_rom[  462] = 'h000007b4; 	    d_addr_rom[  462] = 'h00000ee4; 	    wdata_rom[  462] = 'hf7f74ed9; 	    wvalid_rom[  462] = 0; 
    i_addr_rom[  463] = 'h00000234; 	    d_addr_rom[  463] = 'h0000084c; 	    wdata_rom[  463] = 'h6472b5ca; 	    wvalid_rom[  463] = 1; 
    i_addr_rom[  464] = 'h00000614; 	    d_addr_rom[  464] = 'h00000ac8; 	    wdata_rom[  464] = 'h61fe6cdf; 	    wvalid_rom[  464] = 0; 
    i_addr_rom[  465] = 'h000000ec; 	    d_addr_rom[  465] = 'h00000a30; 	    wdata_rom[  465] = 'h47e09dd6; 	    wvalid_rom[  465] = 1; 
    i_addr_rom[  466] = 'h00000604; 	    d_addr_rom[  466] = 'h00000eb8; 	    wdata_rom[  466] = 'hb0690f43; 	    wvalid_rom[  466] = 0; 
    i_addr_rom[  467] = 'h000006f4; 	    d_addr_rom[  467] = 'h00000ec8; 	    wdata_rom[  467] = 'he3e6b6b9; 	    wvalid_rom[  467] = 1; 
    i_addr_rom[  468] = 'h00000480; 	    d_addr_rom[  468] = 'h00000e00; 	    wdata_rom[  468] = 'h1208c673; 	    wvalid_rom[  468] = 1; 
    i_addr_rom[  469] = 'h00000314; 	    d_addr_rom[  469] = 'h00000a20; 	    wdata_rom[  469] = 'hd5daf357; 	    wvalid_rom[  469] = 0; 
    i_addr_rom[  470] = 'h000007cc; 	    d_addr_rom[  470] = 'h00000d64; 	    wdata_rom[  470] = 'hb1e272d1; 	    wvalid_rom[  470] = 0; 
    i_addr_rom[  471] = 'h00000724; 	    d_addr_rom[  471] = 'h00000dc8; 	    wdata_rom[  471] = 'hbd9701b4; 	    wvalid_rom[  471] = 0; 
    i_addr_rom[  472] = 'h00000444; 	    d_addr_rom[  472] = 'h00000c54; 	    wdata_rom[  472] = 'hcb449066; 	    wvalid_rom[  472] = 1; 
    i_addr_rom[  473] = 'h00000360; 	    d_addr_rom[  473] = 'h00000924; 	    wdata_rom[  473] = 'h6de8dc01; 	    wvalid_rom[  473] = 0; 
    i_addr_rom[  474] = 'h00000018; 	    d_addr_rom[  474] = 'h00000850; 	    wdata_rom[  474] = 'hc5dbe4af; 	    wvalid_rom[  474] = 1; 
    i_addr_rom[  475] = 'h00000278; 	    d_addr_rom[  475] = 'h00000e78; 	    wdata_rom[  475] = 'hba2a0e3c; 	    wvalid_rom[  475] = 0; 
    i_addr_rom[  476] = 'h00000774; 	    d_addr_rom[  476] = 'h00000ae0; 	    wdata_rom[  476] = 'hb29087d8; 	    wvalid_rom[  476] = 0; 
    i_addr_rom[  477] = 'h00000514; 	    d_addr_rom[  477] = 'h00000fe8; 	    wdata_rom[  477] = 'hb480c6f0; 	    wvalid_rom[  477] = 1; 
    i_addr_rom[  478] = 'h00000554; 	    d_addr_rom[  478] = 'h00000f64; 	    wdata_rom[  478] = 'heef70b30; 	    wvalid_rom[  478] = 1; 
    i_addr_rom[  479] = 'h0000043c; 	    d_addr_rom[  479] = 'h00000910; 	    wdata_rom[  479] = 'h8e9b041d; 	    wvalid_rom[  479] = 0; 
    i_addr_rom[  480] = 'h00000764; 	    d_addr_rom[  480] = 'h00000930; 	    wdata_rom[  480] = 'h1b76a018; 	    wvalid_rom[  480] = 0; 
    i_addr_rom[  481] = 'h00000428; 	    d_addr_rom[  481] = 'h00000b28; 	    wdata_rom[  481] = 'hf35e4d6b; 	    wvalid_rom[  481] = 0; 
    i_addr_rom[  482] = 'h000005c4; 	    d_addr_rom[  482] = 'h00000d54; 	    wdata_rom[  482] = 'h2306555e; 	    wvalid_rom[  482] = 0; 
    i_addr_rom[  483] = 'h00000044; 	    d_addr_rom[  483] = 'h00000e90; 	    wdata_rom[  483] = 'h1b29694c; 	    wvalid_rom[  483] = 0; 
    i_addr_rom[  484] = 'h00000314; 	    d_addr_rom[  484] = 'h00000be8; 	    wdata_rom[  484] = 'h03c45310; 	    wvalid_rom[  484] = 1; 
    i_addr_rom[  485] = 'h00000514; 	    d_addr_rom[  485] = 'h00000fd0; 	    wdata_rom[  485] = 'hcac6aace; 	    wvalid_rom[  485] = 1; 
    i_addr_rom[  486] = 'h000003a4; 	    d_addr_rom[  486] = 'h00000a58; 	    wdata_rom[  486] = 'h8d9c2f76; 	    wvalid_rom[  486] = 0; 
    i_addr_rom[  487] = 'h000003ac; 	    d_addr_rom[  487] = 'h00000988; 	    wdata_rom[  487] = 'h1ff24ac6; 	    wvalid_rom[  487] = 0; 
    i_addr_rom[  488] = 'h000004b0; 	    d_addr_rom[  488] = 'h00000bb4; 	    wdata_rom[  488] = 'h4faac0fb; 	    wvalid_rom[  488] = 1; 
    i_addr_rom[  489] = 'h00000484; 	    d_addr_rom[  489] = 'h00000edc; 	    wdata_rom[  489] = 'h62ad4b5b; 	    wvalid_rom[  489] = 1; 
    i_addr_rom[  490] = 'h000001ec; 	    d_addr_rom[  490] = 'h00000a74; 	    wdata_rom[  490] = 'h31a76ca4; 	    wvalid_rom[  490] = 0; 
    i_addr_rom[  491] = 'h000005cc; 	    d_addr_rom[  491] = 'h000009d4; 	    wdata_rom[  491] = 'hf073faea; 	    wvalid_rom[  491] = 1; 
    i_addr_rom[  492] = 'h00000224; 	    d_addr_rom[  492] = 'h000008e0; 	    wdata_rom[  492] = 'he64168fb; 	    wvalid_rom[  492] = 1; 
    i_addr_rom[  493] = 'h00000648; 	    d_addr_rom[  493] = 'h00000c2c; 	    wdata_rom[  493] = 'hd7d55a0e; 	    wvalid_rom[  493] = 0; 
    i_addr_rom[  494] = 'h0000016c; 	    d_addr_rom[  494] = 'h00000b88; 	    wdata_rom[  494] = 'h5522a000; 	    wvalid_rom[  494] = 0; 
    i_addr_rom[  495] = 'h00000218; 	    d_addr_rom[  495] = 'h00000d00; 	    wdata_rom[  495] = 'hfac1164b; 	    wvalid_rom[  495] = 1; 
    i_addr_rom[  496] = 'h000005dc; 	    d_addr_rom[  496] = 'h00000f7c; 	    wdata_rom[  496] = 'h11a16932; 	    wvalid_rom[  496] = 0; 
    i_addr_rom[  497] = 'h0000051c; 	    d_addr_rom[  497] = 'h00000f00; 	    wdata_rom[  497] = 'h126dfcdd; 	    wvalid_rom[  497] = 0; 
    i_addr_rom[  498] = 'h0000037c; 	    d_addr_rom[  498] = 'h00000e6c; 	    wdata_rom[  498] = 'he6fefde5; 	    wvalid_rom[  498] = 0; 
    i_addr_rom[  499] = 'h00000228; 	    d_addr_rom[  499] = 'h00000fa8; 	    wdata_rom[  499] = 'h54aa2115; 	    wvalid_rom[  499] = 1; 
    i_addr_rom[  500] = 'h000003cc; 	    d_addr_rom[  500] = 'h00000db0; 	    wdata_rom[  500] = 'h759b2de2; 	    wvalid_rom[  500] = 0; 
    i_addr_rom[  501] = 'h00000484; 	    d_addr_rom[  501] = 'h00000ae8; 	    wdata_rom[  501] = 'h95c85e02; 	    wvalid_rom[  501] = 0; 
    i_addr_rom[  502] = 'h00000730; 	    d_addr_rom[  502] = 'h00000824; 	    wdata_rom[  502] = 'h066e4e29; 	    wvalid_rom[  502] = 1; 
    i_addr_rom[  503] = 'h00000494; 	    d_addr_rom[  503] = 'h00000af0; 	    wdata_rom[  503] = 'hbc5e06c0; 	    wvalid_rom[  503] = 0; 
    i_addr_rom[  504] = 'h000003e8; 	    d_addr_rom[  504] = 'h00000cd8; 	    wdata_rom[  504] = 'hccf7e426; 	    wvalid_rom[  504] = 1; 
    i_addr_rom[  505] = 'h00000004; 	    d_addr_rom[  505] = 'h00000cb8; 	    wdata_rom[  505] = 'hf3203165; 	    wvalid_rom[  505] = 0; 
    i_addr_rom[  506] = 'h00000578; 	    d_addr_rom[  506] = 'h00000b88; 	    wdata_rom[  506] = 'h1acba77d; 	    wvalid_rom[  506] = 0; 
    i_addr_rom[  507] = 'h000005d0; 	    d_addr_rom[  507] = 'h000008c8; 	    wdata_rom[  507] = 'hefc01f32; 	    wvalid_rom[  507] = 0; 
    i_addr_rom[  508] = 'h00000324; 	    d_addr_rom[  508] = 'h00000ccc; 	    wdata_rom[  508] = 'h57091ff1; 	    wvalid_rom[  508] = 1; 
    i_addr_rom[  509] = 'h00000454; 	    d_addr_rom[  509] = 'h00000b4c; 	    wdata_rom[  509] = 'hcf038504; 	    wvalid_rom[  509] = 0; 
    i_addr_rom[  510] = 'h000003f8; 	    d_addr_rom[  510] = 'h00000a28; 	    wdata_rom[  510] = 'h06dee88a; 	    wvalid_rom[  510] = 0; 
    i_addr_rom[  511] = 'h000003ec; 	    d_addr_rom[  511] = 'h00000c3c; 	    wdata_rom[  511] = 'h9d710ad2; 	    wvalid_rom[  511] = 1; 
    i_addr_rom[  512] = 'h00000160; 	    d_addr_rom[  512] = 'h00000b44; 	    wdata_rom[  512] = 'h6449d5b8; 	    wvalid_rom[  512] = 1; 
    i_addr_rom[  513] = 'h000002c4; 	    d_addr_rom[  513] = 'h00000f44; 	    wdata_rom[  513] = 'hedc96852; 	    wvalid_rom[  513] = 1; 
    i_addr_rom[  514] = 'h00000424; 	    d_addr_rom[  514] = 'h00000ab4; 	    wdata_rom[  514] = 'hb0987a7b; 	    wvalid_rom[  514] = 0; 
    i_addr_rom[  515] = 'h00000258; 	    d_addr_rom[  515] = 'h00000a44; 	    wdata_rom[  515] = 'h3213a8a1; 	    wvalid_rom[  515] = 0; 
    i_addr_rom[  516] = 'h000006e8; 	    d_addr_rom[  516] = 'h00000ab4; 	    wdata_rom[  516] = 'h1e1f26ec; 	    wvalid_rom[  516] = 1; 
    i_addr_rom[  517] = 'h00000278; 	    d_addr_rom[  517] = 'h00000960; 	    wdata_rom[  517] = 'h3345ea2e; 	    wvalid_rom[  517] = 0; 
    i_addr_rom[  518] = 'h000003d8; 	    d_addr_rom[  518] = 'h00000b84; 	    wdata_rom[  518] = 'hc1104109; 	    wvalid_rom[  518] = 1; 
    i_addr_rom[  519] = 'h000005a8; 	    d_addr_rom[  519] = 'h00000b50; 	    wdata_rom[  519] = 'hc4b48aa2; 	    wvalid_rom[  519] = 0; 
    i_addr_rom[  520] = 'h000000cc; 	    d_addr_rom[  520] = 'h00000b24; 	    wdata_rom[  520] = 'ha424a5c8; 	    wvalid_rom[  520] = 1; 
    i_addr_rom[  521] = 'h000005f0; 	    d_addr_rom[  521] = 'h00000d84; 	    wdata_rom[  521] = 'h51c684e7; 	    wvalid_rom[  521] = 0; 
    i_addr_rom[  522] = 'h00000274; 	    d_addr_rom[  522] = 'h000008b8; 	    wdata_rom[  522] = 'hef528fda; 	    wvalid_rom[  522] = 1; 
    i_addr_rom[  523] = 'h00000128; 	    d_addr_rom[  523] = 'h00000d50; 	    wdata_rom[  523] = 'h80df9511; 	    wvalid_rom[  523] = 1; 
    i_addr_rom[  524] = 'h0000038c; 	    d_addr_rom[  524] = 'h00000874; 	    wdata_rom[  524] = 'h1407fb02; 	    wvalid_rom[  524] = 1; 
    i_addr_rom[  525] = 'h000004f0; 	    d_addr_rom[  525] = 'h00000e80; 	    wdata_rom[  525] = 'h4925b1ac; 	    wvalid_rom[  525] = 0; 
    i_addr_rom[  526] = 'h0000061c; 	    d_addr_rom[  526] = 'h00000868; 	    wdata_rom[  526] = 'h3915f208; 	    wvalid_rom[  526] = 1; 
    i_addr_rom[  527] = 'h000007f8; 	    d_addr_rom[  527] = 'h00000d60; 	    wdata_rom[  527] = 'h8af7eecc; 	    wvalid_rom[  527] = 1; 
    i_addr_rom[  528] = 'h000002cc; 	    d_addr_rom[  528] = 'h00000a30; 	    wdata_rom[  528] = 'h14de3a7a; 	    wvalid_rom[  528] = 1; 
    i_addr_rom[  529] = 'h00000090; 	    d_addr_rom[  529] = 'h00000a14; 	    wdata_rom[  529] = 'hefef5712; 	    wvalid_rom[  529] = 1; 
    i_addr_rom[  530] = 'h000004a4; 	    d_addr_rom[  530] = 'h00000b74; 	    wdata_rom[  530] = 'h6b59da49; 	    wvalid_rom[  530] = 1; 
    i_addr_rom[  531] = 'h000006b0; 	    d_addr_rom[  531] = 'h00000d10; 	    wdata_rom[  531] = 'hbb1e432d; 	    wvalid_rom[  531] = 0; 
    i_addr_rom[  532] = 'h0000060c; 	    d_addr_rom[  532] = 'h00000984; 	    wdata_rom[  532] = 'hef70826d; 	    wvalid_rom[  532] = 1; 
    i_addr_rom[  533] = 'h000006b4; 	    d_addr_rom[  533] = 'h00000dfc; 	    wdata_rom[  533] = 'h7d6be8ba; 	    wvalid_rom[  533] = 0; 
    i_addr_rom[  534] = 'h000000f0; 	    d_addr_rom[  534] = 'h000008e4; 	    wdata_rom[  534] = 'hb8bf7fcf; 	    wvalid_rom[  534] = 0; 
    i_addr_rom[  535] = 'h00000308; 	    d_addr_rom[  535] = 'h00000aa0; 	    wdata_rom[  535] = 'hf056b9e9; 	    wvalid_rom[  535] = 0; 
    i_addr_rom[  536] = 'h00000138; 	    d_addr_rom[  536] = 'h00000f98; 	    wdata_rom[  536] = 'h9f20c0d2; 	    wvalid_rom[  536] = 0; 
    i_addr_rom[  537] = 'h00000428; 	    d_addr_rom[  537] = 'h00000e50; 	    wdata_rom[  537] = 'h146cfb49; 	    wvalid_rom[  537] = 1; 
    i_addr_rom[  538] = 'h000006f8; 	    d_addr_rom[  538] = 'h00000888; 	    wdata_rom[  538] = 'hce762b64; 	    wvalid_rom[  538] = 1; 
    i_addr_rom[  539] = 'h000005ac; 	    d_addr_rom[  539] = 'h00000bf0; 	    wdata_rom[  539] = 'h24b1e15c; 	    wvalid_rom[  539] = 1; 
    i_addr_rom[  540] = 'h00000398; 	    d_addr_rom[  540] = 'h000009a4; 	    wdata_rom[  540] = 'h4386c979; 	    wvalid_rom[  540] = 0; 
    i_addr_rom[  541] = 'h00000304; 	    d_addr_rom[  541] = 'h00000cb4; 	    wdata_rom[  541] = 'h649f4efa; 	    wvalid_rom[  541] = 0; 
    i_addr_rom[  542] = 'h00000174; 	    d_addr_rom[  542] = 'h00000838; 	    wdata_rom[  542] = 'h62cb0055; 	    wvalid_rom[  542] = 0; 
    i_addr_rom[  543] = 'h0000016c; 	    d_addr_rom[  543] = 'h00000ff0; 	    wdata_rom[  543] = 'ha252680f; 	    wvalid_rom[  543] = 0; 
    i_addr_rom[  544] = 'h0000035c; 	    d_addr_rom[  544] = 'h00000e8c; 	    wdata_rom[  544] = 'h90135b2c; 	    wvalid_rom[  544] = 1; 
    i_addr_rom[  545] = 'h0000048c; 	    d_addr_rom[  545] = 'h00000d24; 	    wdata_rom[  545] = 'head89aca; 	    wvalid_rom[  545] = 0; 
    i_addr_rom[  546] = 'h000007d0; 	    d_addr_rom[  546] = 'h00000e58; 	    wdata_rom[  546] = 'hbe1bdcca; 	    wvalid_rom[  546] = 1; 
    i_addr_rom[  547] = 'h000004a4; 	    d_addr_rom[  547] = 'h0000096c; 	    wdata_rom[  547] = 'h221b255b; 	    wvalid_rom[  547] = 1; 
    i_addr_rom[  548] = 'h000004d8; 	    d_addr_rom[  548] = 'h00000b90; 	    wdata_rom[  548] = 'hfd5e1468; 	    wvalid_rom[  548] = 0; 
    i_addr_rom[  549] = 'h000001cc; 	    d_addr_rom[  549] = 'h00000f38; 	    wdata_rom[  549] = 'he69664e4; 	    wvalid_rom[  549] = 1; 
    i_addr_rom[  550] = 'h000003b8; 	    d_addr_rom[  550] = 'h00000c10; 	    wdata_rom[  550] = 'hc8a2b8aa; 	    wvalid_rom[  550] = 1; 
    i_addr_rom[  551] = 'h000000ec; 	    d_addr_rom[  551] = 'h000008fc; 	    wdata_rom[  551] = 'haeab6bda; 	    wvalid_rom[  551] = 1; 
    i_addr_rom[  552] = 'h000002d4; 	    d_addr_rom[  552] = 'h000009bc; 	    wdata_rom[  552] = 'hefab45ec; 	    wvalid_rom[  552] = 1; 
    i_addr_rom[  553] = 'h00000450; 	    d_addr_rom[  553] = 'h00000a98; 	    wdata_rom[  553] = 'hf60f5279; 	    wvalid_rom[  553] = 1; 
    i_addr_rom[  554] = 'h0000035c; 	    d_addr_rom[  554] = 'h00000fec; 	    wdata_rom[  554] = 'hf5f54ebf; 	    wvalid_rom[  554] = 1; 
    i_addr_rom[  555] = 'h000001d0; 	    d_addr_rom[  555] = 'h00000a7c; 	    wdata_rom[  555] = 'hac96ccef; 	    wvalid_rom[  555] = 1; 
    i_addr_rom[  556] = 'h000000c4; 	    d_addr_rom[  556] = 'h00000f1c; 	    wdata_rom[  556] = 'h80847fd4; 	    wvalid_rom[  556] = 0; 
    i_addr_rom[  557] = 'h0000003c; 	    d_addr_rom[  557] = 'h00000f2c; 	    wdata_rom[  557] = 'h564a0265; 	    wvalid_rom[  557] = 0; 
    i_addr_rom[  558] = 'h000001c4; 	    d_addr_rom[  558] = 'h00000910; 	    wdata_rom[  558] = 'ha1ac1997; 	    wvalid_rom[  558] = 0; 
    i_addr_rom[  559] = 'h00000514; 	    d_addr_rom[  559] = 'h00000e68; 	    wdata_rom[  559] = 'h32b5d592; 	    wvalid_rom[  559] = 0; 
    i_addr_rom[  560] = 'h00000484; 	    d_addr_rom[  560] = 'h00000bf4; 	    wdata_rom[  560] = 'h6803d59e; 	    wvalid_rom[  560] = 0; 
    i_addr_rom[  561] = 'h000006c8; 	    d_addr_rom[  561] = 'h00000d50; 	    wdata_rom[  561] = 'hc829255e; 	    wvalid_rom[  561] = 1; 
    i_addr_rom[  562] = 'h00000748; 	    d_addr_rom[  562] = 'h000009a8; 	    wdata_rom[  562] = 'hcfa7469a; 	    wvalid_rom[  562] = 0; 
    i_addr_rom[  563] = 'h0000073c; 	    d_addr_rom[  563] = 'h00000b44; 	    wdata_rom[  563] = 'hc517a4b8; 	    wvalid_rom[  563] = 0; 
    i_addr_rom[  564] = 'h000003d0; 	    d_addr_rom[  564] = 'h00000c04; 	    wdata_rom[  564] = 'h66fdadcc; 	    wvalid_rom[  564] = 0; 
    i_addr_rom[  565] = 'h0000043c; 	    d_addr_rom[  565] = 'h000008fc; 	    wdata_rom[  565] = 'hf7b7c234; 	    wvalid_rom[  565] = 1; 
    i_addr_rom[  566] = 'h000007dc; 	    d_addr_rom[  566] = 'h00000f78; 	    wdata_rom[  566] = 'h8cfa424e; 	    wvalid_rom[  566] = 1; 
    i_addr_rom[  567] = 'h0000016c; 	    d_addr_rom[  567] = 'h00000924; 	    wdata_rom[  567] = 'h5288a805; 	    wvalid_rom[  567] = 1; 
    i_addr_rom[  568] = 'h00000704; 	    d_addr_rom[  568] = 'h00000cec; 	    wdata_rom[  568] = 'ha419f950; 	    wvalid_rom[  568] = 0; 
    i_addr_rom[  569] = 'h00000704; 	    d_addr_rom[  569] = 'h00000e78; 	    wdata_rom[  569] = 'hdd54311d; 	    wvalid_rom[  569] = 0; 
    i_addr_rom[  570] = 'h000006c4; 	    d_addr_rom[  570] = 'h00000b5c; 	    wdata_rom[  570] = 'hc36ee4ba; 	    wvalid_rom[  570] = 0; 
    i_addr_rom[  571] = 'h000002b0; 	    d_addr_rom[  571] = 'h00000b78; 	    wdata_rom[  571] = 'h348c5b09; 	    wvalid_rom[  571] = 1; 
    i_addr_rom[  572] = 'h00000600; 	    d_addr_rom[  572] = 'h00000d84; 	    wdata_rom[  572] = 'h8383555f; 	    wvalid_rom[  572] = 1; 
    i_addr_rom[  573] = 'h000000dc; 	    d_addr_rom[  573] = 'h0000091c; 	    wdata_rom[  573] = 'h21b95474; 	    wvalid_rom[  573] = 1; 
    i_addr_rom[  574] = 'h00000484; 	    d_addr_rom[  574] = 'h00000dc8; 	    wdata_rom[  574] = 'he2054bf5; 	    wvalid_rom[  574] = 0; 
    i_addr_rom[  575] = 'h00000204; 	    d_addr_rom[  575] = 'h00000814; 	    wdata_rom[  575] = 'h5b1abdbd; 	    wvalid_rom[  575] = 1; 
    i_addr_rom[  576] = 'h000003a4; 	    d_addr_rom[  576] = 'h00000c68; 	    wdata_rom[  576] = 'hbaac5741; 	    wvalid_rom[  576] = 1; 
    i_addr_rom[  577] = 'h000002b0; 	    d_addr_rom[  577] = 'h00000c5c; 	    wdata_rom[  577] = 'h270248cd; 	    wvalid_rom[  577] = 1; 
    i_addr_rom[  578] = 'h000006c0; 	    d_addr_rom[  578] = 'h00000bd8; 	    wdata_rom[  578] = 'h1babdaf6; 	    wvalid_rom[  578] = 0; 
    i_addr_rom[  579] = 'h000005fc; 	    d_addr_rom[  579] = 'h00000b3c; 	    wdata_rom[  579] = 'hbb2063d0; 	    wvalid_rom[  579] = 1; 
    i_addr_rom[  580] = 'h0000036c; 	    d_addr_rom[  580] = 'h00000f94; 	    wdata_rom[  580] = 'h4b17ca2a; 	    wvalid_rom[  580] = 1; 
    i_addr_rom[  581] = 'h000003f4; 	    d_addr_rom[  581] = 'h00000b98; 	    wdata_rom[  581] = 'h46e8887b; 	    wvalid_rom[  581] = 1; 
    i_addr_rom[  582] = 'h00000310; 	    d_addr_rom[  582] = 'h00000d38; 	    wdata_rom[  582] = 'hab14171c; 	    wvalid_rom[  582] = 0; 
    i_addr_rom[  583] = 'h00000350; 	    d_addr_rom[  583] = 'h00000aa0; 	    wdata_rom[  583] = 'he621e64f; 	    wvalid_rom[  583] = 1; 
    i_addr_rom[  584] = 'h000006cc; 	    d_addr_rom[  584] = 'h00000b20; 	    wdata_rom[  584] = 'h950e38cc; 	    wvalid_rom[  584] = 1; 
    i_addr_rom[  585] = 'h0000059c; 	    d_addr_rom[  585] = 'h00000b38; 	    wdata_rom[  585] = 'h93c030d1; 	    wvalid_rom[  585] = 0; 
    i_addr_rom[  586] = 'h00000188; 	    d_addr_rom[  586] = 'h00000cd0; 	    wdata_rom[  586] = 'hcf17b26f; 	    wvalid_rom[  586] = 0; 
    i_addr_rom[  587] = 'h00000534; 	    d_addr_rom[  587] = 'h00000b98; 	    wdata_rom[  587] = 'h360a0aeb; 	    wvalid_rom[  587] = 0; 
    i_addr_rom[  588] = 'h00000764; 	    d_addr_rom[  588] = 'h00000f70; 	    wdata_rom[  588] = 'h498b0494; 	    wvalid_rom[  588] = 1; 
    i_addr_rom[  589] = 'h00000228; 	    d_addr_rom[  589] = 'h00000838; 	    wdata_rom[  589] = 'hf08679db; 	    wvalid_rom[  589] = 0; 
    i_addr_rom[  590] = 'h000000ec; 	    d_addr_rom[  590] = 'h00000998; 	    wdata_rom[  590] = 'h057e772d; 	    wvalid_rom[  590] = 1; 
    i_addr_rom[  591] = 'h00000468; 	    d_addr_rom[  591] = 'h00000acc; 	    wdata_rom[  591] = 'h5027e293; 	    wvalid_rom[  591] = 0; 
    i_addr_rom[  592] = 'h00000254; 	    d_addr_rom[  592] = 'h00000d60; 	    wdata_rom[  592] = 'h40b1c4e8; 	    wvalid_rom[  592] = 1; 
    i_addr_rom[  593] = 'h0000031c; 	    d_addr_rom[  593] = 'h00000830; 	    wdata_rom[  593] = 'hc2b611a8; 	    wvalid_rom[  593] = 1; 
    i_addr_rom[  594] = 'h00000144; 	    d_addr_rom[  594] = 'h00000f80; 	    wdata_rom[  594] = 'h378b7f7e; 	    wvalid_rom[  594] = 1; 
    i_addr_rom[  595] = 'h000005e0; 	    d_addr_rom[  595] = 'h00000a0c; 	    wdata_rom[  595] = 'h9c5345e4; 	    wvalid_rom[  595] = 0; 
    i_addr_rom[  596] = 'h00000168; 	    d_addr_rom[  596] = 'h00000aec; 	    wdata_rom[  596] = 'h5b26b258; 	    wvalid_rom[  596] = 0; 
    i_addr_rom[  597] = 'h000007d4; 	    d_addr_rom[  597] = 'h00000ff4; 	    wdata_rom[  597] = 'h61169220; 	    wvalid_rom[  597] = 0; 
    i_addr_rom[  598] = 'h00000714; 	    d_addr_rom[  598] = 'h00000ffc; 	    wdata_rom[  598] = 'h9637ae57; 	    wvalid_rom[  598] = 0; 
    i_addr_rom[  599] = 'h00000230; 	    d_addr_rom[  599] = 'h00000b2c; 	    wdata_rom[  599] = 'h6f6b0454; 	    wvalid_rom[  599] = 1; 
    i_addr_rom[  600] = 'h00000238; 	    d_addr_rom[  600] = 'h00000dd8; 	    wdata_rom[  600] = 'h18cfae1d; 	    wvalid_rom[  600] = 1; 
    i_addr_rom[  601] = 'h00000144; 	    d_addr_rom[  601] = 'h00000fd0; 	    wdata_rom[  601] = 'hc2965fe0; 	    wvalid_rom[  601] = 0; 
    i_addr_rom[  602] = 'h0000010c; 	    d_addr_rom[  602] = 'h00000e5c; 	    wdata_rom[  602] = 'hd035e2e0; 	    wvalid_rom[  602] = 0; 
    i_addr_rom[  603] = 'h00000460; 	    d_addr_rom[  603] = 'h00000d6c; 	    wdata_rom[  603] = 'h10b0ef84; 	    wvalid_rom[  603] = 1; 
    i_addr_rom[  604] = 'h000004b8; 	    d_addr_rom[  604] = 'h00000b74; 	    wdata_rom[  604] = 'hc59e5ae1; 	    wvalid_rom[  604] = 0; 
    i_addr_rom[  605] = 'h00000340; 	    d_addr_rom[  605] = 'h00000a58; 	    wdata_rom[  605] = 'h537730cd; 	    wvalid_rom[  605] = 1; 
    i_addr_rom[  606] = 'h00000320; 	    d_addr_rom[  606] = 'h00000994; 	    wdata_rom[  606] = 'h1631ff26; 	    wvalid_rom[  606] = 1; 
    i_addr_rom[  607] = 'h00000344; 	    d_addr_rom[  607] = 'h00000830; 	    wdata_rom[  607] = 'hc1c2d9fa; 	    wvalid_rom[  607] = 1; 
    i_addr_rom[  608] = 'h00000214; 	    d_addr_rom[  608] = 'h00000c98; 	    wdata_rom[  608] = 'h0af1f344; 	    wvalid_rom[  608] = 0; 
    i_addr_rom[  609] = 'h00000780; 	    d_addr_rom[  609] = 'h00000914; 	    wdata_rom[  609] = 'h6d7a36d0; 	    wvalid_rom[  609] = 1; 
    i_addr_rom[  610] = 'h00000670; 	    d_addr_rom[  610] = 'h00000970; 	    wdata_rom[  610] = 'h5511935f; 	    wvalid_rom[  610] = 0; 
    i_addr_rom[  611] = 'h0000055c; 	    d_addr_rom[  611] = 'h000009a4; 	    wdata_rom[  611] = 'hc6b4f7e0; 	    wvalid_rom[  611] = 0; 
    i_addr_rom[  612] = 'h000007c4; 	    d_addr_rom[  612] = 'h00000c00; 	    wdata_rom[  612] = 'h9c943dfd; 	    wvalid_rom[  612] = 0; 
    i_addr_rom[  613] = 'h00000190; 	    d_addr_rom[  613] = 'h00000aec; 	    wdata_rom[  613] = 'hc3e6407c; 	    wvalid_rom[  613] = 1; 
    i_addr_rom[  614] = 'h000000d0; 	    d_addr_rom[  614] = 'h00000df4; 	    wdata_rom[  614] = 'h0f483d4d; 	    wvalid_rom[  614] = 1; 
    i_addr_rom[  615] = 'h00000480; 	    d_addr_rom[  615] = 'h00000988; 	    wdata_rom[  615] = 'h6ee8d9d9; 	    wvalid_rom[  615] = 1; 
    i_addr_rom[  616] = 'h00000324; 	    d_addr_rom[  616] = 'h00000f28; 	    wdata_rom[  616] = 'hac510c28; 	    wvalid_rom[  616] = 1; 
    i_addr_rom[  617] = 'h000001dc; 	    d_addr_rom[  617] = 'h00000cac; 	    wdata_rom[  617] = 'h31c2e94e; 	    wvalid_rom[  617] = 1; 
    i_addr_rom[  618] = 'h000000a0; 	    d_addr_rom[  618] = 'h00000958; 	    wdata_rom[  618] = 'hadc7a2fd; 	    wvalid_rom[  618] = 1; 
    i_addr_rom[  619] = 'h0000029c; 	    d_addr_rom[  619] = 'h00000a40; 	    wdata_rom[  619] = 'h6ce928c2; 	    wvalid_rom[  619] = 0; 
    i_addr_rom[  620] = 'h0000056c; 	    d_addr_rom[  620] = 'h000008cc; 	    wdata_rom[  620] = 'h5efac579; 	    wvalid_rom[  620] = 0; 
    i_addr_rom[  621] = 'h00000074; 	    d_addr_rom[  621] = 'h00000c0c; 	    wdata_rom[  621] = 'hd7a87882; 	    wvalid_rom[  621] = 1; 
    i_addr_rom[  622] = 'h00000008; 	    d_addr_rom[  622] = 'h00000c98; 	    wdata_rom[  622] = 'h9ee610d8; 	    wvalid_rom[  622] = 1; 
    i_addr_rom[  623] = 'h00000230; 	    d_addr_rom[  623] = 'h00000d70; 	    wdata_rom[  623] = 'h33d320ec; 	    wvalid_rom[  623] = 1; 
    i_addr_rom[  624] = 'h000005b4; 	    d_addr_rom[  624] = 'h00000bc4; 	    wdata_rom[  624] = 'heba499e2; 	    wvalid_rom[  624] = 1; 
    i_addr_rom[  625] = 'h00000658; 	    d_addr_rom[  625] = 'h000009ac; 	    wdata_rom[  625] = 'hda1eaf4a; 	    wvalid_rom[  625] = 1; 
    i_addr_rom[  626] = 'h000006bc; 	    d_addr_rom[  626] = 'h000008c0; 	    wdata_rom[  626] = 'h70390cb1; 	    wvalid_rom[  626] = 1; 
    i_addr_rom[  627] = 'h00000178; 	    d_addr_rom[  627] = 'h00000c88; 	    wdata_rom[  627] = 'h32cc46fe; 	    wvalid_rom[  627] = 1; 
    i_addr_rom[  628] = 'h00000694; 	    d_addr_rom[  628] = 'h00000d8c; 	    wdata_rom[  628] = 'h757bf011; 	    wvalid_rom[  628] = 1; 
    i_addr_rom[  629] = 'h000002b4; 	    d_addr_rom[  629] = 'h00000d04; 	    wdata_rom[  629] = 'h272ab5c4; 	    wvalid_rom[  629] = 0; 
    i_addr_rom[  630] = 'h00000320; 	    d_addr_rom[  630] = 'h00000888; 	    wdata_rom[  630] = 'h4e05a1ad; 	    wvalid_rom[  630] = 0; 
    i_addr_rom[  631] = 'h000006ac; 	    d_addr_rom[  631] = 'h00000f98; 	    wdata_rom[  631] = 'h31933bd2; 	    wvalid_rom[  631] = 0; 
    i_addr_rom[  632] = 'h00000154; 	    d_addr_rom[  632] = 'h00000fe4; 	    wdata_rom[  632] = 'hc19539c8; 	    wvalid_rom[  632] = 1; 
    i_addr_rom[  633] = 'h000002a0; 	    d_addr_rom[  633] = 'h00000a84; 	    wdata_rom[  633] = 'h7c945ede; 	    wvalid_rom[  633] = 0; 
    i_addr_rom[  634] = 'h00000588; 	    d_addr_rom[  634] = 'h00000ba0; 	    wdata_rom[  634] = 'hbeb5bb4f; 	    wvalid_rom[  634] = 1; 
    i_addr_rom[  635] = 'h000007b8; 	    d_addr_rom[  635] = 'h00000dcc; 	    wdata_rom[  635] = 'haf7a74d8; 	    wvalid_rom[  635] = 0; 
    i_addr_rom[  636] = 'h000003dc; 	    d_addr_rom[  636] = 'h00000f54; 	    wdata_rom[  636] = 'h0b3e8846; 	    wvalid_rom[  636] = 0; 
    i_addr_rom[  637] = 'h00000390; 	    d_addr_rom[  637] = 'h00000e50; 	    wdata_rom[  637] = 'h61198811; 	    wvalid_rom[  637] = 1; 
    i_addr_rom[  638] = 'h00000528; 	    d_addr_rom[  638] = 'h00000d70; 	    wdata_rom[  638] = 'hd6769a6a; 	    wvalid_rom[  638] = 1; 
    i_addr_rom[  639] = 'h000000e8; 	    d_addr_rom[  639] = 'h00000c30; 	    wdata_rom[  639] = 'h85aa059d; 	    wvalid_rom[  639] = 1; 
    i_addr_rom[  640] = 'h000004e4; 	    d_addr_rom[  640] = 'h00000e94; 	    wdata_rom[  640] = 'h1a09aa51; 	    wvalid_rom[  640] = 1; 
    i_addr_rom[  641] = 'h00000158; 	    d_addr_rom[  641] = 'h00000f74; 	    wdata_rom[  641] = 'h518203f2; 	    wvalid_rom[  641] = 0; 
    i_addr_rom[  642] = 'h000003cc; 	    d_addr_rom[  642] = 'h00000de0; 	    wdata_rom[  642] = 'h82885cf8; 	    wvalid_rom[  642] = 1; 
    i_addr_rom[  643] = 'h000006c0; 	    d_addr_rom[  643] = 'h00000c2c; 	    wdata_rom[  643] = 'h52d2aef3; 	    wvalid_rom[  643] = 1; 
    i_addr_rom[  644] = 'h000007e0; 	    d_addr_rom[  644] = 'h00000a34; 	    wdata_rom[  644] = 'h28c3b066; 	    wvalid_rom[  644] = 0; 
    i_addr_rom[  645] = 'h00000438; 	    d_addr_rom[  645] = 'h00000a7c; 	    wdata_rom[  645] = 'h0fbe024c; 	    wvalid_rom[  645] = 1; 
    i_addr_rom[  646] = 'h00000268; 	    d_addr_rom[  646] = 'h00000fbc; 	    wdata_rom[  646] = 'h28fb41c2; 	    wvalid_rom[  646] = 0; 
    i_addr_rom[  647] = 'h0000043c; 	    d_addr_rom[  647] = 'h00000d24; 	    wdata_rom[  647] = 'h6851cb68; 	    wvalid_rom[  647] = 0; 
    i_addr_rom[  648] = 'h000005c0; 	    d_addr_rom[  648] = 'h00000d88; 	    wdata_rom[  648] = 'h1783c0f3; 	    wvalid_rom[  648] = 1; 
    i_addr_rom[  649] = 'h000003e0; 	    d_addr_rom[  649] = 'h00000b84; 	    wdata_rom[  649] = 'h7d5c464a; 	    wvalid_rom[  649] = 0; 
    i_addr_rom[  650] = 'h000003b0; 	    d_addr_rom[  650] = 'h00000f34; 	    wdata_rom[  650] = 'hc3ede311; 	    wvalid_rom[  650] = 0; 
    i_addr_rom[  651] = 'h000001ec; 	    d_addr_rom[  651] = 'h00000dcc; 	    wdata_rom[  651] = 'h5f81368f; 	    wvalid_rom[  651] = 0; 
    i_addr_rom[  652] = 'h000004f0; 	    d_addr_rom[  652] = 'h00000838; 	    wdata_rom[  652] = 'h27aa075d; 	    wvalid_rom[  652] = 0; 
    i_addr_rom[  653] = 'h00000354; 	    d_addr_rom[  653] = 'h00000b80; 	    wdata_rom[  653] = 'ha418dab6; 	    wvalid_rom[  653] = 0; 
    i_addr_rom[  654] = 'h00000694; 	    d_addr_rom[  654] = 'h00000804; 	    wdata_rom[  654] = 'hd5673445; 	    wvalid_rom[  654] = 0; 
    i_addr_rom[  655] = 'h0000013c; 	    d_addr_rom[  655] = 'h00000d6c; 	    wdata_rom[  655] = 'hac522bb3; 	    wvalid_rom[  655] = 0; 
    i_addr_rom[  656] = 'h00000624; 	    d_addr_rom[  656] = 'h000008b4; 	    wdata_rom[  656] = 'h9bbaf41d; 	    wvalid_rom[  656] = 0; 
    i_addr_rom[  657] = 'h00000700; 	    d_addr_rom[  657] = 'h00000820; 	    wdata_rom[  657] = 'h1782a40d; 	    wvalid_rom[  657] = 0; 
    i_addr_rom[  658] = 'h00000588; 	    d_addr_rom[  658] = 'h000009a0; 	    wdata_rom[  658] = 'h421130bf; 	    wvalid_rom[  658] = 1; 
    i_addr_rom[  659] = 'h0000030c; 	    d_addr_rom[  659] = 'h00000b54; 	    wdata_rom[  659] = 'hc3faca54; 	    wvalid_rom[  659] = 1; 
    i_addr_rom[  660] = 'h00000604; 	    d_addr_rom[  660] = 'h00000dc4; 	    wdata_rom[  660] = 'hf6209b1e; 	    wvalid_rom[  660] = 1; 
    i_addr_rom[  661] = 'h000002a0; 	    d_addr_rom[  661] = 'h00000fe4; 	    wdata_rom[  661] = 'h6599ddc2; 	    wvalid_rom[  661] = 1; 
    i_addr_rom[  662] = 'h000006f4; 	    d_addr_rom[  662] = 'h00000abc; 	    wdata_rom[  662] = 'h31a09250; 	    wvalid_rom[  662] = 0; 
    i_addr_rom[  663] = 'h000002cc; 	    d_addr_rom[  663] = 'h000008f8; 	    wdata_rom[  663] = 'h35b53c55; 	    wvalid_rom[  663] = 0; 
    i_addr_rom[  664] = 'h00000618; 	    d_addr_rom[  664] = 'h00000b84; 	    wdata_rom[  664] = 'hbf3a02cc; 	    wvalid_rom[  664] = 1; 
    i_addr_rom[  665] = 'h000007c8; 	    d_addr_rom[  665] = 'h00000c80; 	    wdata_rom[  665] = 'h733bdda2; 	    wvalid_rom[  665] = 0; 
    i_addr_rom[  666] = 'h000007d0; 	    d_addr_rom[  666] = 'h00000e68; 	    wdata_rom[  666] = 'h634132f2; 	    wvalid_rom[  666] = 0; 
    i_addr_rom[  667] = 'h000007cc; 	    d_addr_rom[  667] = 'h00000d38; 	    wdata_rom[  667] = 'h712cbb19; 	    wvalid_rom[  667] = 1; 
    i_addr_rom[  668] = 'h00000784; 	    d_addr_rom[  668] = 'h00000e84; 	    wdata_rom[  668] = 'hccd36744; 	    wvalid_rom[  668] = 0; 
    i_addr_rom[  669] = 'h00000480; 	    d_addr_rom[  669] = 'h00000920; 	    wdata_rom[  669] = 'h94401b98; 	    wvalid_rom[  669] = 0; 
    i_addr_rom[  670] = 'h0000053c; 	    d_addr_rom[  670] = 'h00000c5c; 	    wdata_rom[  670] = 'he819752a; 	    wvalid_rom[  670] = 0; 
    i_addr_rom[  671] = 'h0000007c; 	    d_addr_rom[  671] = 'h00000b48; 	    wdata_rom[  671] = 'h6d7fa785; 	    wvalid_rom[  671] = 1; 
    i_addr_rom[  672] = 'h000001e8; 	    d_addr_rom[  672] = 'h00000848; 	    wdata_rom[  672] = 'h1e0dbd8f; 	    wvalid_rom[  672] = 0; 
    i_addr_rom[  673] = 'h00000684; 	    d_addr_rom[  673] = 'h00000e50; 	    wdata_rom[  673] = 'hac6be192; 	    wvalid_rom[  673] = 1; 
    i_addr_rom[  674] = 'h00000064; 	    d_addr_rom[  674] = 'h00000a1c; 	    wdata_rom[  674] = 'h23296b07; 	    wvalid_rom[  674] = 0; 
    i_addr_rom[  675] = 'h00000574; 	    d_addr_rom[  675] = 'h00000910; 	    wdata_rom[  675] = 'h21abf494; 	    wvalid_rom[  675] = 0; 
    i_addr_rom[  676] = 'h0000026c; 	    d_addr_rom[  676] = 'h00000ae0; 	    wdata_rom[  676] = 'ha3d532e0; 	    wvalid_rom[  676] = 0; 
    i_addr_rom[  677] = 'h000000b0; 	    d_addr_rom[  677] = 'h00000a80; 	    wdata_rom[  677] = 'hbbde8d4f; 	    wvalid_rom[  677] = 1; 
    i_addr_rom[  678] = 'h000006c8; 	    d_addr_rom[  678] = 'h00000838; 	    wdata_rom[  678] = 'hc1afc16e; 	    wvalid_rom[  678] = 1; 
    i_addr_rom[  679] = 'h000003a4; 	    d_addr_rom[  679] = 'h00000904; 	    wdata_rom[  679] = 'h103e25be; 	    wvalid_rom[  679] = 0; 
    i_addr_rom[  680] = 'h00000164; 	    d_addr_rom[  680] = 'h00000e98; 	    wdata_rom[  680] = 'hc39b1ca9; 	    wvalid_rom[  680] = 0; 
    i_addr_rom[  681] = 'h0000005c; 	    d_addr_rom[  681] = 'h00000eb4; 	    wdata_rom[  681] = 'h94d4011e; 	    wvalid_rom[  681] = 1; 
    i_addr_rom[  682] = 'h00000110; 	    d_addr_rom[  682] = 'h00000ff0; 	    wdata_rom[  682] = 'h60e5aec3; 	    wvalid_rom[  682] = 1; 
    i_addr_rom[  683] = 'h000005c0; 	    d_addr_rom[  683] = 'h00000d14; 	    wdata_rom[  683] = 'hfb5398ba; 	    wvalid_rom[  683] = 0; 
    i_addr_rom[  684] = 'h000006e8; 	    d_addr_rom[  684] = 'h00000b8c; 	    wdata_rom[  684] = 'hc2508bb7; 	    wvalid_rom[  684] = 1; 
    i_addr_rom[  685] = 'h000007d4; 	    d_addr_rom[  685] = 'h00000994; 	    wdata_rom[  685] = 'h0099efa1; 	    wvalid_rom[  685] = 1; 
    i_addr_rom[  686] = 'h000005f8; 	    d_addr_rom[  686] = 'h00000840; 	    wdata_rom[  686] = 'hb339232a; 	    wvalid_rom[  686] = 0; 
    i_addr_rom[  687] = 'h000001cc; 	    d_addr_rom[  687] = 'h00000fc4; 	    wdata_rom[  687] = 'haea46e36; 	    wvalid_rom[  687] = 0; 
    i_addr_rom[  688] = 'h000005a4; 	    d_addr_rom[  688] = 'h000009fc; 	    wdata_rom[  688] = 'h02f1460d; 	    wvalid_rom[  688] = 0; 
    i_addr_rom[  689] = 'h0000065c; 	    d_addr_rom[  689] = 'h00000b00; 	    wdata_rom[  689] = 'hc28d5a7b; 	    wvalid_rom[  689] = 0; 
    i_addr_rom[  690] = 'h000007c8; 	    d_addr_rom[  690] = 'h00000e44; 	    wdata_rom[  690] = 'hb013c70a; 	    wvalid_rom[  690] = 0; 
    i_addr_rom[  691] = 'h0000033c; 	    d_addr_rom[  691] = 'h000009a0; 	    wdata_rom[  691] = 'h40e29ce5; 	    wvalid_rom[  691] = 0; 
    i_addr_rom[  692] = 'h000007b8; 	    d_addr_rom[  692] = 'h00000cb8; 	    wdata_rom[  692] = 'hcefd9434; 	    wvalid_rom[  692] = 1; 
    i_addr_rom[  693] = 'h00000368; 	    d_addr_rom[  693] = 'h00000b24; 	    wdata_rom[  693] = 'ha1cd8cdb; 	    wvalid_rom[  693] = 1; 
    i_addr_rom[  694] = 'h000002f8; 	    d_addr_rom[  694] = 'h00000d58; 	    wdata_rom[  694] = 'h67fcad97; 	    wvalid_rom[  694] = 0; 
    i_addr_rom[  695] = 'h0000059c; 	    d_addr_rom[  695] = 'h00000d7c; 	    wdata_rom[  695] = 'h9cacdb74; 	    wvalid_rom[  695] = 0; 
    i_addr_rom[  696] = 'h0000067c; 	    d_addr_rom[  696] = 'h00000e24; 	    wdata_rom[  696] = 'h10e01f0d; 	    wvalid_rom[  696] = 0; 
    i_addr_rom[  697] = 'h000004e4; 	    d_addr_rom[  697] = 'h00000940; 	    wdata_rom[  697] = 'h0a32e90f; 	    wvalid_rom[  697] = 1; 
    i_addr_rom[  698] = 'h000003b8; 	    d_addr_rom[  698] = 'h00000810; 	    wdata_rom[  698] = 'h700ff2ae; 	    wvalid_rom[  698] = 0; 
    i_addr_rom[  699] = 'h00000220; 	    d_addr_rom[  699] = 'h00000dac; 	    wdata_rom[  699] = 'h373a68ed; 	    wvalid_rom[  699] = 1; 
    i_addr_rom[  700] = 'h0000062c; 	    d_addr_rom[  700] = 'h00000890; 	    wdata_rom[  700] = 'h65677bee; 	    wvalid_rom[  700] = 1; 
    i_addr_rom[  701] = 'h0000033c; 	    d_addr_rom[  701] = 'h00000bcc; 	    wdata_rom[  701] = 'h35564d1e; 	    wvalid_rom[  701] = 1; 
    i_addr_rom[  702] = 'h000004ac; 	    d_addr_rom[  702] = 'h00000a7c; 	    wdata_rom[  702] = 'hb0c80469; 	    wvalid_rom[  702] = 1; 
    i_addr_rom[  703] = 'h00000694; 	    d_addr_rom[  703] = 'h00000c30; 	    wdata_rom[  703] = 'hdce6bd55; 	    wvalid_rom[  703] = 1; 
    i_addr_rom[  704] = 'h0000036c; 	    d_addr_rom[  704] = 'h000009a8; 	    wdata_rom[  704] = 'h939f96be; 	    wvalid_rom[  704] = 0; 
    i_addr_rom[  705] = 'h00000350; 	    d_addr_rom[  705] = 'h00000bd4; 	    wdata_rom[  705] = 'hd95b2ed3; 	    wvalid_rom[  705] = 1; 
    i_addr_rom[  706] = 'h00000348; 	    d_addr_rom[  706] = 'h00000dd4; 	    wdata_rom[  706] = 'h6b03b9b9; 	    wvalid_rom[  706] = 0; 
    i_addr_rom[  707] = 'h000004b0; 	    d_addr_rom[  707] = 'h00000cd0; 	    wdata_rom[  707] = 'h81b3ddc5; 	    wvalid_rom[  707] = 0; 
    i_addr_rom[  708] = 'h00000744; 	    d_addr_rom[  708] = 'h00000a84; 	    wdata_rom[  708] = 'hfc4eff6a; 	    wvalid_rom[  708] = 0; 
    i_addr_rom[  709] = 'h00000330; 	    d_addr_rom[  709] = 'h00000cc0; 	    wdata_rom[  709] = 'h47a01d3e; 	    wvalid_rom[  709] = 0; 
    i_addr_rom[  710] = 'h00000668; 	    d_addr_rom[  710] = 'h00000fa8; 	    wdata_rom[  710] = 'he9af4951; 	    wvalid_rom[  710] = 0; 
    i_addr_rom[  711] = 'h000002b4; 	    d_addr_rom[  711] = 'h00000f44; 	    wdata_rom[  711] = 'h8bae2f4f; 	    wvalid_rom[  711] = 1; 
    i_addr_rom[  712] = 'h00000768; 	    d_addr_rom[  712] = 'h00000998; 	    wdata_rom[  712] = 'h39a83672; 	    wvalid_rom[  712] = 1; 
    i_addr_rom[  713] = 'h00000028; 	    d_addr_rom[  713] = 'h00000c3c; 	    wdata_rom[  713] = 'h7ed213af; 	    wvalid_rom[  713] = 1; 
    i_addr_rom[  714] = 'h000000e4; 	    d_addr_rom[  714] = 'h00000f24; 	    wdata_rom[  714] = 'hdaa6e297; 	    wvalid_rom[  714] = 0; 
    i_addr_rom[  715] = 'h00000580; 	    d_addr_rom[  715] = 'h00000d50; 	    wdata_rom[  715] = 'h7fc2da96; 	    wvalid_rom[  715] = 0; 
    i_addr_rom[  716] = 'h00000374; 	    d_addr_rom[  716] = 'h00000b94; 	    wdata_rom[  716] = 'h0abe131e; 	    wvalid_rom[  716] = 1; 
    i_addr_rom[  717] = 'h000007a0; 	    d_addr_rom[  717] = 'h00000e90; 	    wdata_rom[  717] = 'h5d17c717; 	    wvalid_rom[  717] = 0; 
    i_addr_rom[  718] = 'h00000454; 	    d_addr_rom[  718] = 'h00000a14; 	    wdata_rom[  718] = 'hbb5c223f; 	    wvalid_rom[  718] = 1; 
    i_addr_rom[  719] = 'h00000660; 	    d_addr_rom[  719] = 'h00000a18; 	    wdata_rom[  719] = 'ha7aa65f5; 	    wvalid_rom[  719] = 0; 
    i_addr_rom[  720] = 'h000005f0; 	    d_addr_rom[  720] = 'h00000870; 	    wdata_rom[  720] = 'h6d1d91e2; 	    wvalid_rom[  720] = 1; 
    i_addr_rom[  721] = 'h000002f4; 	    d_addr_rom[  721] = 'h00000da8; 	    wdata_rom[  721] = 'h3b42a8ce; 	    wvalid_rom[  721] = 0; 
    i_addr_rom[  722] = 'h00000798; 	    d_addr_rom[  722] = 'h00000b54; 	    wdata_rom[  722] = 'ha68a1df4; 	    wvalid_rom[  722] = 1; 
    i_addr_rom[  723] = 'h00000068; 	    d_addr_rom[  723] = 'h00000c48; 	    wdata_rom[  723] = 'h7deafcec; 	    wvalid_rom[  723] = 0; 
    i_addr_rom[  724] = 'h0000056c; 	    d_addr_rom[  724] = 'h00000a7c; 	    wdata_rom[  724] = 'h5b094ba3; 	    wvalid_rom[  724] = 0; 
    i_addr_rom[  725] = 'h00000178; 	    d_addr_rom[  725] = 'h00000db4; 	    wdata_rom[  725] = 'h548c4098; 	    wvalid_rom[  725] = 1; 
    i_addr_rom[  726] = 'h00000580; 	    d_addr_rom[  726] = 'h0000086c; 	    wdata_rom[  726] = 'h571ccaa4; 	    wvalid_rom[  726] = 0; 
    i_addr_rom[  727] = 'h00000154; 	    d_addr_rom[  727] = 'h00000c60; 	    wdata_rom[  727] = 'h5ab2db64; 	    wvalid_rom[  727] = 0; 
    i_addr_rom[  728] = 'h000000a0; 	    d_addr_rom[  728] = 'h00000f0c; 	    wdata_rom[  728] = 'hcb997bfa; 	    wvalid_rom[  728] = 1; 
    i_addr_rom[  729] = 'h00000368; 	    d_addr_rom[  729] = 'h0000082c; 	    wdata_rom[  729] = 'haad8d803; 	    wvalid_rom[  729] = 1; 
    i_addr_rom[  730] = 'h00000474; 	    d_addr_rom[  730] = 'h00000c34; 	    wdata_rom[  730] = 'h27d37af8; 	    wvalid_rom[  730] = 1; 
    i_addr_rom[  731] = 'h000007dc; 	    d_addr_rom[  731] = 'h000008a4; 	    wdata_rom[  731] = 'ha13a8450; 	    wvalid_rom[  731] = 1; 
    i_addr_rom[  732] = 'h000001bc; 	    d_addr_rom[  732] = 'h00000cb4; 	    wdata_rom[  732] = 'h7dd5571a; 	    wvalid_rom[  732] = 1; 
    i_addr_rom[  733] = 'h000007dc; 	    d_addr_rom[  733] = 'h000008d4; 	    wdata_rom[  733] = 'h2b038680; 	    wvalid_rom[  733] = 1; 
    i_addr_rom[  734] = 'h000005dc; 	    d_addr_rom[  734] = 'h00000c30; 	    wdata_rom[  734] = 'h3bb0b32b; 	    wvalid_rom[  734] = 1; 
    i_addr_rom[  735] = 'h000001fc; 	    d_addr_rom[  735] = 'h00000a14; 	    wdata_rom[  735] = 'h9c173d74; 	    wvalid_rom[  735] = 0; 
    i_addr_rom[  736] = 'h0000077c; 	    d_addr_rom[  736] = 'h00000d68; 	    wdata_rom[  736] = 'h28fe02e3; 	    wvalid_rom[  736] = 1; 
    i_addr_rom[  737] = 'h00000294; 	    d_addr_rom[  737] = 'h00000fe0; 	    wdata_rom[  737] = 'h5389188e; 	    wvalid_rom[  737] = 0; 
    i_addr_rom[  738] = 'h00000384; 	    d_addr_rom[  738] = 'h0000085c; 	    wdata_rom[  738] = 'h4b38157b; 	    wvalid_rom[  738] = 0; 
    i_addr_rom[  739] = 'h000002cc; 	    d_addr_rom[  739] = 'h00000cd0; 	    wdata_rom[  739] = 'h30725c66; 	    wvalid_rom[  739] = 0; 
    i_addr_rom[  740] = 'h00000280; 	    d_addr_rom[  740] = 'h00000908; 	    wdata_rom[  740] = 'hb9541b33; 	    wvalid_rom[  740] = 1; 
    i_addr_rom[  741] = 'h000005a8; 	    d_addr_rom[  741] = 'h00000dfc; 	    wdata_rom[  741] = 'h7fffa388; 	    wvalid_rom[  741] = 1; 
    i_addr_rom[  742] = 'h00000694; 	    d_addr_rom[  742] = 'h00000b5c; 	    wdata_rom[  742] = 'h533387c9; 	    wvalid_rom[  742] = 0; 
    i_addr_rom[  743] = 'h00000238; 	    d_addr_rom[  743] = 'h00000ff8; 	    wdata_rom[  743] = 'h3a3600f3; 	    wvalid_rom[  743] = 1; 
    i_addr_rom[  744] = 'h000002e0; 	    d_addr_rom[  744] = 'h00000b60; 	    wdata_rom[  744] = 'h83157c07; 	    wvalid_rom[  744] = 1; 
    i_addr_rom[  745] = 'h00000640; 	    d_addr_rom[  745] = 'h00000adc; 	    wdata_rom[  745] = 'h2f6c4216; 	    wvalid_rom[  745] = 1; 
    i_addr_rom[  746] = 'h0000065c; 	    d_addr_rom[  746] = 'h00000850; 	    wdata_rom[  746] = 'hda695fa7; 	    wvalid_rom[  746] = 0; 
    i_addr_rom[  747] = 'h0000066c; 	    d_addr_rom[  747] = 'h00000e94; 	    wdata_rom[  747] = 'h610dabe4; 	    wvalid_rom[  747] = 0; 
    i_addr_rom[  748] = 'h0000075c; 	    d_addr_rom[  748] = 'h00000c40; 	    wdata_rom[  748] = 'hb70936a0; 	    wvalid_rom[  748] = 1; 
    i_addr_rom[  749] = 'h000000fc; 	    d_addr_rom[  749] = 'h00000cdc; 	    wdata_rom[  749] = 'h3f949dea; 	    wvalid_rom[  749] = 0; 
    i_addr_rom[  750] = 'h00000600; 	    d_addr_rom[  750] = 'h00000850; 	    wdata_rom[  750] = 'hcf19461c; 	    wvalid_rom[  750] = 0; 
    i_addr_rom[  751] = 'h0000041c; 	    d_addr_rom[  751] = 'h00000d7c; 	    wdata_rom[  751] = 'ha9881585; 	    wvalid_rom[  751] = 0; 
    i_addr_rom[  752] = 'h0000045c; 	    d_addr_rom[  752] = 'h00000f88; 	    wdata_rom[  752] = 'ha12dcac5; 	    wvalid_rom[  752] = 1; 
    i_addr_rom[  753] = 'h00000330; 	    d_addr_rom[  753] = 'h00000b30; 	    wdata_rom[  753] = 'h7d4cd427; 	    wvalid_rom[  753] = 0; 
    i_addr_rom[  754] = 'h00000048; 	    d_addr_rom[  754] = 'h00000bbc; 	    wdata_rom[  754] = 'h0a327e52; 	    wvalid_rom[  754] = 0; 
    i_addr_rom[  755] = 'h000002b8; 	    d_addr_rom[  755] = 'h00000ecc; 	    wdata_rom[  755] = 'hfd44d9d6; 	    wvalid_rom[  755] = 1; 
    i_addr_rom[  756] = 'h000006c0; 	    d_addr_rom[  756] = 'h00000954; 	    wdata_rom[  756] = 'h30dbc00f; 	    wvalid_rom[  756] = 1; 
    i_addr_rom[  757] = 'h00000610; 	    d_addr_rom[  757] = 'h00000f38; 	    wdata_rom[  757] = 'h21921b29; 	    wvalid_rom[  757] = 1; 
    i_addr_rom[  758] = 'h000007c0; 	    d_addr_rom[  758] = 'h00000d18; 	    wdata_rom[  758] = 'h5eef2bda; 	    wvalid_rom[  758] = 1; 
    i_addr_rom[  759] = 'h0000043c; 	    d_addr_rom[  759] = 'h00000fec; 	    wdata_rom[  759] = 'hda34d0c9; 	    wvalid_rom[  759] = 1; 
    i_addr_rom[  760] = 'h00000008; 	    d_addr_rom[  760] = 'h00000adc; 	    wdata_rom[  760] = 'h6bfa4479; 	    wvalid_rom[  760] = 1; 
    i_addr_rom[  761] = 'h0000063c; 	    d_addr_rom[  761] = 'h00000ff4; 	    wdata_rom[  761] = 'hd3cbf815; 	    wvalid_rom[  761] = 1; 
    i_addr_rom[  762] = 'h00000018; 	    d_addr_rom[  762] = 'h00000d44; 	    wdata_rom[  762] = 'h951a257d; 	    wvalid_rom[  762] = 1; 
    i_addr_rom[  763] = 'h000003a4; 	    d_addr_rom[  763] = 'h00000ab4; 	    wdata_rom[  763] = 'hcc3f1862; 	    wvalid_rom[  763] = 0; 
    i_addr_rom[  764] = 'h00000514; 	    d_addr_rom[  764] = 'h000009d4; 	    wdata_rom[  764] = 'h32127c98; 	    wvalid_rom[  764] = 1; 
    i_addr_rom[  765] = 'h000003b0; 	    d_addr_rom[  765] = 'h00000b6c; 	    wdata_rom[  765] = 'hc847c68c; 	    wvalid_rom[  765] = 0; 
    i_addr_rom[  766] = 'h000006c0; 	    d_addr_rom[  766] = 'h00000ae8; 	    wdata_rom[  766] = 'h52da06a5; 	    wvalid_rom[  766] = 0; 
    i_addr_rom[  767] = 'h000004c8; 	    d_addr_rom[  767] = 'h00000f80; 	    wdata_rom[  767] = 'hd50de680; 	    wvalid_rom[  767] = 1; 
    i_addr_rom[  768] = 'h000006d4; 	    d_addr_rom[  768] = 'h00000df0; 	    wdata_rom[  768] = 'hf6213d0f; 	    wvalid_rom[  768] = 0; 
    i_addr_rom[  769] = 'h0000062c; 	    d_addr_rom[  769] = 'h00000ab0; 	    wdata_rom[  769] = 'h77ebb822; 	    wvalid_rom[  769] = 0; 
    i_addr_rom[  770] = 'h000007b0; 	    d_addr_rom[  770] = 'h00000c64; 	    wdata_rom[  770] = 'h679a267e; 	    wvalid_rom[  770] = 1; 
    i_addr_rom[  771] = 'h00000200; 	    d_addr_rom[  771] = 'h0000097c; 	    wdata_rom[  771] = 'h6700862d; 	    wvalid_rom[  771] = 1; 
    i_addr_rom[  772] = 'h00000118; 	    d_addr_rom[  772] = 'h00000c64; 	    wdata_rom[  772] = 'h8746dedb; 	    wvalid_rom[  772] = 0; 
    i_addr_rom[  773] = 'h00000390; 	    d_addr_rom[  773] = 'h000009b0; 	    wdata_rom[  773] = 'h1a86adf3; 	    wvalid_rom[  773] = 1; 
    i_addr_rom[  774] = 'h0000068c; 	    d_addr_rom[  774] = 'h00000874; 	    wdata_rom[  774] = 'hee0ae711; 	    wvalid_rom[  774] = 1; 
    i_addr_rom[  775] = 'h00000224; 	    d_addr_rom[  775] = 'h00000874; 	    wdata_rom[  775] = 'hbe866f36; 	    wvalid_rom[  775] = 1; 
    i_addr_rom[  776] = 'h000002cc; 	    d_addr_rom[  776] = 'h0000096c; 	    wdata_rom[  776] = 'hd01abbc3; 	    wvalid_rom[  776] = 1; 
    i_addr_rom[  777] = 'h0000003c; 	    d_addr_rom[  777] = 'h00000ce4; 	    wdata_rom[  777] = 'h6b91983c; 	    wvalid_rom[  777] = 1; 
    i_addr_rom[  778] = 'h00000094; 	    d_addr_rom[  778] = 'h00000e04; 	    wdata_rom[  778] = 'h03449dae; 	    wvalid_rom[  778] = 0; 
    i_addr_rom[  779] = 'h000003a8; 	    d_addr_rom[  779] = 'h00000a04; 	    wdata_rom[  779] = 'hf44c1c40; 	    wvalid_rom[  779] = 1; 
    i_addr_rom[  780] = 'h00000420; 	    d_addr_rom[  780] = 'h00000d9c; 	    wdata_rom[  780] = 'h3fdcfff4; 	    wvalid_rom[  780] = 0; 
    i_addr_rom[  781] = 'h000005f0; 	    d_addr_rom[  781] = 'h0000097c; 	    wdata_rom[  781] = 'hdb6436bb; 	    wvalid_rom[  781] = 0; 
    i_addr_rom[  782] = 'h00000578; 	    d_addr_rom[  782] = 'h00000c4c; 	    wdata_rom[  782] = 'hbe1ac80d; 	    wvalid_rom[  782] = 1; 
    i_addr_rom[  783] = 'h000000f0; 	    d_addr_rom[  783] = 'h000009b4; 	    wdata_rom[  783] = 'h6a1c58bd; 	    wvalid_rom[  783] = 1; 
    i_addr_rom[  784] = 'h00000738; 	    d_addr_rom[  784] = 'h00000dc8; 	    wdata_rom[  784] = 'h13fb717e; 	    wvalid_rom[  784] = 0; 
    i_addr_rom[  785] = 'h000000a8; 	    d_addr_rom[  785] = 'h00000d3c; 	    wdata_rom[  785] = 'h524a1bbe; 	    wvalid_rom[  785] = 1; 
    i_addr_rom[  786] = 'h00000270; 	    d_addr_rom[  786] = 'h00000954; 	    wdata_rom[  786] = 'h13ca3704; 	    wvalid_rom[  786] = 0; 
    i_addr_rom[  787] = 'h000000fc; 	    d_addr_rom[  787] = 'h00000aa8; 	    wdata_rom[  787] = 'hc2c6adb4; 	    wvalid_rom[  787] = 0; 
    i_addr_rom[  788] = 'h0000002c; 	    d_addr_rom[  788] = 'h00000898; 	    wdata_rom[  788] = 'hf933518c; 	    wvalid_rom[  788] = 0; 
    i_addr_rom[  789] = 'h00000364; 	    d_addr_rom[  789] = 'h00000bfc; 	    wdata_rom[  789] = 'h88609d22; 	    wvalid_rom[  789] = 0; 
    i_addr_rom[  790] = 'h00000128; 	    d_addr_rom[  790] = 'h00000d18; 	    wdata_rom[  790] = 'he629d762; 	    wvalid_rom[  790] = 0; 
    i_addr_rom[  791] = 'h000006ec; 	    d_addr_rom[  791] = 'h00000a68; 	    wdata_rom[  791] = 'h53ddef75; 	    wvalid_rom[  791] = 0; 
    i_addr_rom[  792] = 'h000006ec; 	    d_addr_rom[  792] = 'h00000b10; 	    wdata_rom[  792] = 'h29190e9c; 	    wvalid_rom[  792] = 1; 
    i_addr_rom[  793] = 'h00000254; 	    d_addr_rom[  793] = 'h00000a40; 	    wdata_rom[  793] = 'h11d1abf9; 	    wvalid_rom[  793] = 1; 
    i_addr_rom[  794] = 'h000001e4; 	    d_addr_rom[  794] = 'h00000b0c; 	    wdata_rom[  794] = 'h3c488543; 	    wvalid_rom[  794] = 1; 
    i_addr_rom[  795] = 'h000006b4; 	    d_addr_rom[  795] = 'h00000bdc; 	    wdata_rom[  795] = 'hfbcc2fb7; 	    wvalid_rom[  795] = 0; 
    i_addr_rom[  796] = 'h000000ac; 	    d_addr_rom[  796] = 'h00000ccc; 	    wdata_rom[  796] = 'h7a5628de; 	    wvalid_rom[  796] = 1; 
    i_addr_rom[  797] = 'h00000508; 	    d_addr_rom[  797] = 'h00000e2c; 	    wdata_rom[  797] = 'he9178211; 	    wvalid_rom[  797] = 0; 
    i_addr_rom[  798] = 'h000002f0; 	    d_addr_rom[  798] = 'h00000b2c; 	    wdata_rom[  798] = 'h8b4d1753; 	    wvalid_rom[  798] = 0; 
    i_addr_rom[  799] = 'h00000768; 	    d_addr_rom[  799] = 'h00000b74; 	    wdata_rom[  799] = 'hfb640a21; 	    wvalid_rom[  799] = 1; 
    i_addr_rom[  800] = 'h00000418; 	    d_addr_rom[  800] = 'h0000096c; 	    wdata_rom[  800] = 'h36f47c94; 	    wvalid_rom[  800] = 0; 
    i_addr_rom[  801] = 'h00000608; 	    d_addr_rom[  801] = 'h00000da4; 	    wdata_rom[  801] = 'hb43ab45b; 	    wvalid_rom[  801] = 1; 
    i_addr_rom[  802] = 'h00000700; 	    d_addr_rom[  802] = 'h00000bcc; 	    wdata_rom[  802] = 'h3449b8e7; 	    wvalid_rom[  802] = 1; 
    i_addr_rom[  803] = 'h0000023c; 	    d_addr_rom[  803] = 'h00000a78; 	    wdata_rom[  803] = 'h4b0c104d; 	    wvalid_rom[  803] = 0; 
    i_addr_rom[  804] = 'h00000360; 	    d_addr_rom[  804] = 'h00000e50; 	    wdata_rom[  804] = 'h8031af95; 	    wvalid_rom[  804] = 1; 
    i_addr_rom[  805] = 'h000000a0; 	    d_addr_rom[  805] = 'h00000a14; 	    wdata_rom[  805] = 'h64d05168; 	    wvalid_rom[  805] = 0; 
    i_addr_rom[  806] = 'h000000f4; 	    d_addr_rom[  806] = 'h00000a30; 	    wdata_rom[  806] = 'h5a4a9989; 	    wvalid_rom[  806] = 0; 
    i_addr_rom[  807] = 'h000006b0; 	    d_addr_rom[  807] = 'h00000e60; 	    wdata_rom[  807] = 'h4853e8df; 	    wvalid_rom[  807] = 0; 
    i_addr_rom[  808] = 'h0000005c; 	    d_addr_rom[  808] = 'h00000a68; 	    wdata_rom[  808] = 'h08ab7af5; 	    wvalid_rom[  808] = 0; 
    i_addr_rom[  809] = 'h00000294; 	    d_addr_rom[  809] = 'h00000b7c; 	    wdata_rom[  809] = 'h66a5464e; 	    wvalid_rom[  809] = 1; 
    i_addr_rom[  810] = 'h000007c4; 	    d_addr_rom[  810] = 'h00000eb8; 	    wdata_rom[  810] = 'hdc0de603; 	    wvalid_rom[  810] = 0; 
    i_addr_rom[  811] = 'h000000b4; 	    d_addr_rom[  811] = 'h00000d24; 	    wdata_rom[  811] = 'h2eaea86b; 	    wvalid_rom[  811] = 0; 
    i_addr_rom[  812] = 'h000007e0; 	    d_addr_rom[  812] = 'h00000da0; 	    wdata_rom[  812] = 'h6f4aeda0; 	    wvalid_rom[  812] = 0; 
    i_addr_rom[  813] = 'h0000077c; 	    d_addr_rom[  813] = 'h00000994; 	    wdata_rom[  813] = 'hcf8f16e1; 	    wvalid_rom[  813] = 1; 
    i_addr_rom[  814] = 'h0000075c; 	    d_addr_rom[  814] = 'h00000b78; 	    wdata_rom[  814] = 'hb0d7dc99; 	    wvalid_rom[  814] = 1; 
    i_addr_rom[  815] = 'h000002d4; 	    d_addr_rom[  815] = 'h00000ab0; 	    wdata_rom[  815] = 'hf0a3f3ff; 	    wvalid_rom[  815] = 0; 
    i_addr_rom[  816] = 'h00000674; 	    d_addr_rom[  816] = 'h00000e58; 	    wdata_rom[  816] = 'h252c2df8; 	    wvalid_rom[  816] = 0; 
    i_addr_rom[  817] = 'h00000340; 	    d_addr_rom[  817] = 'h00000cc4; 	    wdata_rom[  817] = 'hb616cf91; 	    wvalid_rom[  817] = 0; 
    i_addr_rom[  818] = 'h00000298; 	    d_addr_rom[  818] = 'h00000e7c; 	    wdata_rom[  818] = 'h57740f2a; 	    wvalid_rom[  818] = 0; 
    i_addr_rom[  819] = 'h00000020; 	    d_addr_rom[  819] = 'h00000b10; 	    wdata_rom[  819] = 'h1b304714; 	    wvalid_rom[  819] = 0; 
    i_addr_rom[  820] = 'h00000520; 	    d_addr_rom[  820] = 'h00000948; 	    wdata_rom[  820] = 'h4f65abec; 	    wvalid_rom[  820] = 0; 
    i_addr_rom[  821] = 'h0000026c; 	    d_addr_rom[  821] = 'h0000087c; 	    wdata_rom[  821] = 'hda2fe8be; 	    wvalid_rom[  821] = 1; 
    i_addr_rom[  822] = 'h00000048; 	    d_addr_rom[  822] = 'h00000e54; 	    wdata_rom[  822] = 'h6907c237; 	    wvalid_rom[  822] = 1; 
    i_addr_rom[  823] = 'h00000564; 	    d_addr_rom[  823] = 'h000009e8; 	    wdata_rom[  823] = 'h50ba7488; 	    wvalid_rom[  823] = 1; 
    i_addr_rom[  824] = 'h00000628; 	    d_addr_rom[  824] = 'h00000b84; 	    wdata_rom[  824] = 'h3703f0d5; 	    wvalid_rom[  824] = 1; 
    i_addr_rom[  825] = 'h00000534; 	    d_addr_rom[  825] = 'h00000f70; 	    wdata_rom[  825] = 'hbff988f7; 	    wvalid_rom[  825] = 1; 
    i_addr_rom[  826] = 'h00000518; 	    d_addr_rom[  826] = 'h00000eb4; 	    wdata_rom[  826] = 'h4d4e5db1; 	    wvalid_rom[  826] = 1; 
    i_addr_rom[  827] = 'h0000009c; 	    d_addr_rom[  827] = 'h00000d2c; 	    wdata_rom[  827] = 'h41ead6bb; 	    wvalid_rom[  827] = 1; 
    i_addr_rom[  828] = 'h00000658; 	    d_addr_rom[  828] = 'h00000ee0; 	    wdata_rom[  828] = 'he6db867f; 	    wvalid_rom[  828] = 0; 
    i_addr_rom[  829] = 'h00000084; 	    d_addr_rom[  829] = 'h00000a7c; 	    wdata_rom[  829] = 'h6bba95c4; 	    wvalid_rom[  829] = 1; 
    i_addr_rom[  830] = 'h00000438; 	    d_addr_rom[  830] = 'h00000e34; 	    wdata_rom[  830] = 'h68c419a6; 	    wvalid_rom[  830] = 0; 
    i_addr_rom[  831] = 'h00000720; 	    d_addr_rom[  831] = 'h00000fd4; 	    wdata_rom[  831] = 'h6c45f25b; 	    wvalid_rom[  831] = 1; 
    i_addr_rom[  832] = 'h0000003c; 	    d_addr_rom[  832] = 'h00000f28; 	    wdata_rom[  832] = 'h436d1def; 	    wvalid_rom[  832] = 1; 
    i_addr_rom[  833] = 'h000003f0; 	    d_addr_rom[  833] = 'h00000bd8; 	    wdata_rom[  833] = 'h06c1c0af; 	    wvalid_rom[  833] = 0; 
    i_addr_rom[  834] = 'h00000510; 	    d_addr_rom[  834] = 'h00000b3c; 	    wdata_rom[  834] = 'h276b1768; 	    wvalid_rom[  834] = 0; 
    i_addr_rom[  835] = 'h00000134; 	    d_addr_rom[  835] = 'h00000fa4; 	    wdata_rom[  835] = 'h87107847; 	    wvalid_rom[  835] = 0; 
    i_addr_rom[  836] = 'h00000014; 	    d_addr_rom[  836] = 'h00000a38; 	    wdata_rom[  836] = 'hb369486c; 	    wvalid_rom[  836] = 0; 
    i_addr_rom[  837] = 'h00000074; 	    d_addr_rom[  837] = 'h00000a54; 	    wdata_rom[  837] = 'h2494009c; 	    wvalid_rom[  837] = 0; 
    i_addr_rom[  838] = 'h00000664; 	    d_addr_rom[  838] = 'h0000080c; 	    wdata_rom[  838] = 'h4f1e30de; 	    wvalid_rom[  838] = 1; 
    i_addr_rom[  839] = 'h000000e0; 	    d_addr_rom[  839] = 'h00000d0c; 	    wdata_rom[  839] = 'hdffea1d1; 	    wvalid_rom[  839] = 0; 
    i_addr_rom[  840] = 'h0000032c; 	    d_addr_rom[  840] = 'h00000afc; 	    wdata_rom[  840] = 'heb785178; 	    wvalid_rom[  840] = 1; 
    i_addr_rom[  841] = 'h000001c0; 	    d_addr_rom[  841] = 'h00000bc0; 	    wdata_rom[  841] = 'hb0801ea5; 	    wvalid_rom[  841] = 1; 
    i_addr_rom[  842] = 'h000003f4; 	    d_addr_rom[  842] = 'h00000918; 	    wdata_rom[  842] = 'hbee85117; 	    wvalid_rom[  842] = 0; 
    i_addr_rom[  843] = 'h00000770; 	    d_addr_rom[  843] = 'h00000ab0; 	    wdata_rom[  843] = 'h692a1fb6; 	    wvalid_rom[  843] = 1; 
    i_addr_rom[  844] = 'h00000550; 	    d_addr_rom[  844] = 'h00000ccc; 	    wdata_rom[  844] = 'hd2493aed; 	    wvalid_rom[  844] = 0; 
    i_addr_rom[  845] = 'h00000424; 	    d_addr_rom[  845] = 'h00000a44; 	    wdata_rom[  845] = 'h97d2c929; 	    wvalid_rom[  845] = 0; 
    i_addr_rom[  846] = 'h00000790; 	    d_addr_rom[  846] = 'h00000f24; 	    wdata_rom[  846] = 'hcd431c24; 	    wvalid_rom[  846] = 0; 
    i_addr_rom[  847] = 'h00000190; 	    d_addr_rom[  847] = 'h00000858; 	    wdata_rom[  847] = 'hc0fba0ad; 	    wvalid_rom[  847] = 1; 
    i_addr_rom[  848] = 'h0000006c; 	    d_addr_rom[  848] = 'h00000f18; 	    wdata_rom[  848] = 'hc8ec01e5; 	    wvalid_rom[  848] = 1; 
    i_addr_rom[  849] = 'h0000040c; 	    d_addr_rom[  849] = 'h00000b9c; 	    wdata_rom[  849] = 'h8266d848; 	    wvalid_rom[  849] = 0; 
    i_addr_rom[  850] = 'h00000670; 	    d_addr_rom[  850] = 'h00000de8; 	    wdata_rom[  850] = 'h66d4d40c; 	    wvalid_rom[  850] = 1; 
    i_addr_rom[  851] = 'h000000c0; 	    d_addr_rom[  851] = 'h00000c04; 	    wdata_rom[  851] = 'h2671771a; 	    wvalid_rom[  851] = 1; 
    i_addr_rom[  852] = 'h00000600; 	    d_addr_rom[  852] = 'h00000b6c; 	    wdata_rom[  852] = 'h6eecec24; 	    wvalid_rom[  852] = 1; 
    i_addr_rom[  853] = 'h0000010c; 	    d_addr_rom[  853] = 'h00000d40; 	    wdata_rom[  853] = 'h1602cd8c; 	    wvalid_rom[  853] = 1; 
    i_addr_rom[  854] = 'h0000005c; 	    d_addr_rom[  854] = 'h00000aa8; 	    wdata_rom[  854] = 'h4859560a; 	    wvalid_rom[  854] = 1; 
    i_addr_rom[  855] = 'h00000560; 	    d_addr_rom[  855] = 'h00000d48; 	    wdata_rom[  855] = 'h7ea39a19; 	    wvalid_rom[  855] = 1; 
    i_addr_rom[  856] = 'h000002e8; 	    d_addr_rom[  856] = 'h00000834; 	    wdata_rom[  856] = 'ha1dd4d40; 	    wvalid_rom[  856] = 0; 
    i_addr_rom[  857] = 'h00000410; 	    d_addr_rom[  857] = 'h00000e20; 	    wdata_rom[  857] = 'hc603c893; 	    wvalid_rom[  857] = 1; 
    i_addr_rom[  858] = 'h0000075c; 	    d_addr_rom[  858] = 'h00000fd0; 	    wdata_rom[  858] = 'hfc21a54d; 	    wvalid_rom[  858] = 0; 
    i_addr_rom[  859] = 'h000005c8; 	    d_addr_rom[  859] = 'h00000fa8; 	    wdata_rom[  859] = 'h7a34a109; 	    wvalid_rom[  859] = 0; 
    i_addr_rom[  860] = 'h00000254; 	    d_addr_rom[  860] = 'h00000ae4; 	    wdata_rom[  860] = 'he0c1d08b; 	    wvalid_rom[  860] = 0; 
    i_addr_rom[  861] = 'h000005e4; 	    d_addr_rom[  861] = 'h000009b4; 	    wdata_rom[  861] = 'heda8e7b0; 	    wvalid_rom[  861] = 0; 
    i_addr_rom[  862] = 'h00000174; 	    d_addr_rom[  862] = 'h00000e80; 	    wdata_rom[  862] = 'h1650b83c; 	    wvalid_rom[  862] = 0; 
    i_addr_rom[  863] = 'h00000598; 	    d_addr_rom[  863] = 'h00000cdc; 	    wdata_rom[  863] = 'hcb025663; 	    wvalid_rom[  863] = 0; 
    i_addr_rom[  864] = 'h000003b4; 	    d_addr_rom[  864] = 'h00000ecc; 	    wdata_rom[  864] = 'h60548499; 	    wvalid_rom[  864] = 1; 
    i_addr_rom[  865] = 'h00000324; 	    d_addr_rom[  865] = 'h00000aac; 	    wdata_rom[  865] = 'h51f95b53; 	    wvalid_rom[  865] = 1; 
    i_addr_rom[  866] = 'h0000014c; 	    d_addr_rom[  866] = 'h00000eb4; 	    wdata_rom[  866] = 'hd8878025; 	    wvalid_rom[  866] = 0; 
    i_addr_rom[  867] = 'h000001d8; 	    d_addr_rom[  867] = 'h00000cb4; 	    wdata_rom[  867] = 'hee7cc6dc; 	    wvalid_rom[  867] = 0; 
    i_addr_rom[  868] = 'h000006a0; 	    d_addr_rom[  868] = 'h0000091c; 	    wdata_rom[  868] = 'hf2ab3409; 	    wvalid_rom[  868] = 1; 
    i_addr_rom[  869] = 'h000001dc; 	    d_addr_rom[  869] = 'h00000818; 	    wdata_rom[  869] = 'h01b13665; 	    wvalid_rom[  869] = 0; 
    i_addr_rom[  870] = 'h000003ac; 	    d_addr_rom[  870] = 'h00000ab8; 	    wdata_rom[  870] = 'h8af3c2d7; 	    wvalid_rom[  870] = 1; 
    i_addr_rom[  871] = 'h00000084; 	    d_addr_rom[  871] = 'h000009cc; 	    wdata_rom[  871] = 'h4db6db91; 	    wvalid_rom[  871] = 0; 
    i_addr_rom[  872] = 'h00000298; 	    d_addr_rom[  872] = 'h00000e40; 	    wdata_rom[  872] = 'hc5c80001; 	    wvalid_rom[  872] = 0; 
    i_addr_rom[  873] = 'h00000788; 	    d_addr_rom[  873] = 'h00000eb8; 	    wdata_rom[  873] = 'he3247abd; 	    wvalid_rom[  873] = 0; 
    i_addr_rom[  874] = 'h000001b8; 	    d_addr_rom[  874] = 'h00000d3c; 	    wdata_rom[  874] = 'hf1dc07f7; 	    wvalid_rom[  874] = 0; 
    i_addr_rom[  875] = 'h00000370; 	    d_addr_rom[  875] = 'h0000082c; 	    wdata_rom[  875] = 'hc590f1bd; 	    wvalid_rom[  875] = 1; 
    i_addr_rom[  876] = 'h00000510; 	    d_addr_rom[  876] = 'h00000de8; 	    wdata_rom[  876] = 'h0cafbd17; 	    wvalid_rom[  876] = 1; 
    i_addr_rom[  877] = 'h000002c4; 	    d_addr_rom[  877] = 'h00000b34; 	    wdata_rom[  877] = 'h380f485b; 	    wvalid_rom[  877] = 1; 
    i_addr_rom[  878] = 'h000005d4; 	    d_addr_rom[  878] = 'h00000984; 	    wdata_rom[  878] = 'ha7ecc584; 	    wvalid_rom[  878] = 1; 
    i_addr_rom[  879] = 'h000006a0; 	    d_addr_rom[  879] = 'h000008a0; 	    wdata_rom[  879] = 'h1805f8fe; 	    wvalid_rom[  879] = 0; 
    i_addr_rom[  880] = 'h00000434; 	    d_addr_rom[  880] = 'h000009c0; 	    wdata_rom[  880] = 'h13ceb57b; 	    wvalid_rom[  880] = 1; 
    i_addr_rom[  881] = 'h00000048; 	    d_addr_rom[  881] = 'h00000d58; 	    wdata_rom[  881] = 'hf038b3de; 	    wvalid_rom[  881] = 0; 
    i_addr_rom[  882] = 'h000003e0; 	    d_addr_rom[  882] = 'h00000a6c; 	    wdata_rom[  882] = 'he936d806; 	    wvalid_rom[  882] = 1; 
    i_addr_rom[  883] = 'h0000000c; 	    d_addr_rom[  883] = 'h00000bb0; 	    wdata_rom[  883] = 'h9f04823c; 	    wvalid_rom[  883] = 1; 
    i_addr_rom[  884] = 'h00000754; 	    d_addr_rom[  884] = 'h00000a94; 	    wdata_rom[  884] = 'hc1ad5436; 	    wvalid_rom[  884] = 0; 
    i_addr_rom[  885] = 'h00000300; 	    d_addr_rom[  885] = 'h00000d48; 	    wdata_rom[  885] = 'hecb4815f; 	    wvalid_rom[  885] = 0; 
    i_addr_rom[  886] = 'h000005dc; 	    d_addr_rom[  886] = 'h00000a8c; 	    wdata_rom[  886] = 'hfecaed14; 	    wvalid_rom[  886] = 0; 
    i_addr_rom[  887] = 'h0000022c; 	    d_addr_rom[  887] = 'h00000800; 	    wdata_rom[  887] = 'h88067858; 	    wvalid_rom[  887] = 1; 
    i_addr_rom[  888] = 'h000001fc; 	    d_addr_rom[  888] = 'h00000ddc; 	    wdata_rom[  888] = 'h03ffdba0; 	    wvalid_rom[  888] = 1; 
    i_addr_rom[  889] = 'h000007a4; 	    d_addr_rom[  889] = 'h00000b2c; 	    wdata_rom[  889] = 'h7af1ec2e; 	    wvalid_rom[  889] = 0; 
    i_addr_rom[  890] = 'h0000030c; 	    d_addr_rom[  890] = 'h00000f2c; 	    wdata_rom[  890] = 'h60c76004; 	    wvalid_rom[  890] = 1; 
    i_addr_rom[  891] = 'h00000538; 	    d_addr_rom[  891] = 'h00000b1c; 	    wdata_rom[  891] = 'h336b70c2; 	    wvalid_rom[  891] = 1; 
    i_addr_rom[  892] = 'h000001f0; 	    d_addr_rom[  892] = 'h00000b78; 	    wdata_rom[  892] = 'hf7465eec; 	    wvalid_rom[  892] = 1; 
    i_addr_rom[  893] = 'h0000046c; 	    d_addr_rom[  893] = 'h000008b4; 	    wdata_rom[  893] = 'h62cc2211; 	    wvalid_rom[  893] = 0; 
    i_addr_rom[  894] = 'h000002a8; 	    d_addr_rom[  894] = 'h00000840; 	    wdata_rom[  894] = 'h0cd2c60b; 	    wvalid_rom[  894] = 0; 
    i_addr_rom[  895] = 'h00000454; 	    d_addr_rom[  895] = 'h00000aa4; 	    wdata_rom[  895] = 'h9fdd7957; 	    wvalid_rom[  895] = 1; 
    i_addr_rom[  896] = 'h00000268; 	    d_addr_rom[  896] = 'h000009c4; 	    wdata_rom[  896] = 'he2b49eb8; 	    wvalid_rom[  896] = 0; 
    i_addr_rom[  897] = 'h00000478; 	    d_addr_rom[  897] = 'h00000c78; 	    wdata_rom[  897] = 'h807fd657; 	    wvalid_rom[  897] = 0; 
    i_addr_rom[  898] = 'h000006a4; 	    d_addr_rom[  898] = 'h00000ef4; 	    wdata_rom[  898] = 'h570cfa86; 	    wvalid_rom[  898] = 1; 
    i_addr_rom[  899] = 'h0000034c; 	    d_addr_rom[  899] = 'h00000f00; 	    wdata_rom[  899] = 'h0bbf62e1; 	    wvalid_rom[  899] = 1; 
    i_addr_rom[  900] = 'h0000030c; 	    d_addr_rom[  900] = 'h00000edc; 	    wdata_rom[  900] = 'hbf7c684f; 	    wvalid_rom[  900] = 1; 
    i_addr_rom[  901] = 'h000002b0; 	    d_addr_rom[  901] = 'h00000a24; 	    wdata_rom[  901] = 'h2365f817; 	    wvalid_rom[  901] = 1; 
    i_addr_rom[  902] = 'h000001a0; 	    d_addr_rom[  902] = 'h00000fbc; 	    wdata_rom[  902] = 'h10089061; 	    wvalid_rom[  902] = 1; 
    i_addr_rom[  903] = 'h000007fc; 	    d_addr_rom[  903] = 'h00000cb8; 	    wdata_rom[  903] = 'hab5e8913; 	    wvalid_rom[  903] = 1; 
    i_addr_rom[  904] = 'h00000608; 	    d_addr_rom[  904] = 'h000009f4; 	    wdata_rom[  904] = 'hba9d7949; 	    wvalid_rom[  904] = 1; 
    i_addr_rom[  905] = 'h00000090; 	    d_addr_rom[  905] = 'h00000c10; 	    wdata_rom[  905] = 'hf1d1b707; 	    wvalid_rom[  905] = 1; 
    i_addr_rom[  906] = 'h00000128; 	    d_addr_rom[  906] = 'h00000d70; 	    wdata_rom[  906] = 'h6ba970e4; 	    wvalid_rom[  906] = 0; 
    i_addr_rom[  907] = 'h00000614; 	    d_addr_rom[  907] = 'h00000fbc; 	    wdata_rom[  907] = 'h85da27cb; 	    wvalid_rom[  907] = 1; 
    i_addr_rom[  908] = 'h0000076c; 	    d_addr_rom[  908] = 'h00000dd8; 	    wdata_rom[  908] = 'hbaefbbd6; 	    wvalid_rom[  908] = 0; 
    i_addr_rom[  909] = 'h00000404; 	    d_addr_rom[  909] = 'h00000bc0; 	    wdata_rom[  909] = 'h024a61ec; 	    wvalid_rom[  909] = 0; 
    i_addr_rom[  910] = 'h000001b8; 	    d_addr_rom[  910] = 'h000008a0; 	    wdata_rom[  910] = 'h2b60b4ec; 	    wvalid_rom[  910] = 1; 
    i_addr_rom[  911] = 'h0000039c; 	    d_addr_rom[  911] = 'h00000ee8; 	    wdata_rom[  911] = 'ha24d85ce; 	    wvalid_rom[  911] = 0; 
    i_addr_rom[  912] = 'h00000778; 	    d_addr_rom[  912] = 'h00000df0; 	    wdata_rom[  912] = 'h464ed375; 	    wvalid_rom[  912] = 1; 
    i_addr_rom[  913] = 'h00000244; 	    d_addr_rom[  913] = 'h00000900; 	    wdata_rom[  913] = 'h98766c08; 	    wvalid_rom[  913] = 1; 
    i_addr_rom[  914] = 'h00000714; 	    d_addr_rom[  914] = 'h00000a78; 	    wdata_rom[  914] = 'hf1f0107c; 	    wvalid_rom[  914] = 1; 
    i_addr_rom[  915] = 'h000001e4; 	    d_addr_rom[  915] = 'h00000a58; 	    wdata_rom[  915] = 'ha340bd95; 	    wvalid_rom[  915] = 0; 
    i_addr_rom[  916] = 'h0000020c; 	    d_addr_rom[  916] = 'h00000b64; 	    wdata_rom[  916] = 'h35455c9f; 	    wvalid_rom[  916] = 0; 
    i_addr_rom[  917] = 'h00000668; 	    d_addr_rom[  917] = 'h000008d4; 	    wdata_rom[  917] = 'hfcd5d9aa; 	    wvalid_rom[  917] = 0; 
    i_addr_rom[  918] = 'h00000298; 	    d_addr_rom[  918] = 'h00000c1c; 	    wdata_rom[  918] = 'h1302ac46; 	    wvalid_rom[  918] = 0; 
    i_addr_rom[  919] = 'h0000024c; 	    d_addr_rom[  919] = 'h0000085c; 	    wdata_rom[  919] = 'hd8de1f39; 	    wvalid_rom[  919] = 1; 
    i_addr_rom[  920] = 'h00000134; 	    d_addr_rom[  920] = 'h00000f94; 	    wdata_rom[  920] = 'h670c056c; 	    wvalid_rom[  920] = 0; 
    i_addr_rom[  921] = 'h00000378; 	    d_addr_rom[  921] = 'h00000854; 	    wdata_rom[  921] = 'hbac4e4de; 	    wvalid_rom[  921] = 0; 
    i_addr_rom[  922] = 'h0000043c; 	    d_addr_rom[  922] = 'h00000abc; 	    wdata_rom[  922] = 'ha498d15e; 	    wvalid_rom[  922] = 1; 
    i_addr_rom[  923] = 'h00000264; 	    d_addr_rom[  923] = 'h00000b64; 	    wdata_rom[  923] = 'h7f7d73b9; 	    wvalid_rom[  923] = 0; 
    i_addr_rom[  924] = 'h000004c0; 	    d_addr_rom[  924] = 'h00000bc8; 	    wdata_rom[  924] = 'hc1d10c7b; 	    wvalid_rom[  924] = 0; 
    i_addr_rom[  925] = 'h000004b8; 	    d_addr_rom[  925] = 'h00000860; 	    wdata_rom[  925] = 'ha1290973; 	    wvalid_rom[  925] = 1; 
    i_addr_rom[  926] = 'h000001b0; 	    d_addr_rom[  926] = 'h00000944; 	    wdata_rom[  926] = 'h443f069c; 	    wvalid_rom[  926] = 0; 
    i_addr_rom[  927] = 'h000007c0; 	    d_addr_rom[  927] = 'h00000b94; 	    wdata_rom[  927] = 'h94e6d139; 	    wvalid_rom[  927] = 0; 
    i_addr_rom[  928] = 'h000005c8; 	    d_addr_rom[  928] = 'h00000930; 	    wdata_rom[  928] = 'h8dcb1b32; 	    wvalid_rom[  928] = 1; 
    i_addr_rom[  929] = 'h00000224; 	    d_addr_rom[  929] = 'h00000e98; 	    wdata_rom[  929] = 'hde8dc275; 	    wvalid_rom[  929] = 0; 
    i_addr_rom[  930] = 'h000007e0; 	    d_addr_rom[  930] = 'h00000848; 	    wdata_rom[  930] = 'hc9ca7c39; 	    wvalid_rom[  930] = 0; 
    i_addr_rom[  931] = 'h00000444; 	    d_addr_rom[  931] = 'h00000e30; 	    wdata_rom[  931] = 'h9efb0c93; 	    wvalid_rom[  931] = 0; 
    i_addr_rom[  932] = 'h00000304; 	    d_addr_rom[  932] = 'h00000f10; 	    wdata_rom[  932] = 'h373cee32; 	    wvalid_rom[  932] = 0; 
    i_addr_rom[  933] = 'h0000023c; 	    d_addr_rom[  933] = 'h00000e34; 	    wdata_rom[  933] = 'h2cb8a2ba; 	    wvalid_rom[  933] = 1; 
    i_addr_rom[  934] = 'h000001fc; 	    d_addr_rom[  934] = 'h00000c48; 	    wdata_rom[  934] = 'h7889ef27; 	    wvalid_rom[  934] = 1; 
    i_addr_rom[  935] = 'h000006f0; 	    d_addr_rom[  935] = 'h00000b18; 	    wdata_rom[  935] = 'hafcd0929; 	    wvalid_rom[  935] = 0; 
    i_addr_rom[  936] = 'h00000438; 	    d_addr_rom[  936] = 'h00000b8c; 	    wdata_rom[  936] = 'h8e7d1432; 	    wvalid_rom[  936] = 0; 
    i_addr_rom[  937] = 'h000001d8; 	    d_addr_rom[  937] = 'h00000d38; 	    wdata_rom[  937] = 'hfbd80f53; 	    wvalid_rom[  937] = 1; 
    i_addr_rom[  938] = 'h00000048; 	    d_addr_rom[  938] = 'h00000bfc; 	    wdata_rom[  938] = 'hc85a4313; 	    wvalid_rom[  938] = 0; 
    i_addr_rom[  939] = 'h00000678; 	    d_addr_rom[  939] = 'h00000840; 	    wdata_rom[  939] = 'heb22fc63; 	    wvalid_rom[  939] = 0; 
    i_addr_rom[  940] = 'h000002e4; 	    d_addr_rom[  940] = 'h00000fc4; 	    wdata_rom[  940] = 'hb21a15bd; 	    wvalid_rom[  940] = 1; 
    i_addr_rom[  941] = 'h00000254; 	    d_addr_rom[  941] = 'h00000a20; 	    wdata_rom[  941] = 'h15c355e6; 	    wvalid_rom[  941] = 1; 
    i_addr_rom[  942] = 'h000000e4; 	    d_addr_rom[  942] = 'h00000920; 	    wdata_rom[  942] = 'haa938572; 	    wvalid_rom[  942] = 0; 
    i_addr_rom[  943] = 'h00000468; 	    d_addr_rom[  943] = 'h00000a48; 	    wdata_rom[  943] = 'hfd4706c4; 	    wvalid_rom[  943] = 1; 
    i_addr_rom[  944] = 'h00000408; 	    d_addr_rom[  944] = 'h00000864; 	    wdata_rom[  944] = 'hd32840f2; 	    wvalid_rom[  944] = 1; 
    i_addr_rom[  945] = 'h000000ac; 	    d_addr_rom[  945] = 'h00000cac; 	    wdata_rom[  945] = 'h8514cc62; 	    wvalid_rom[  945] = 1; 
    i_addr_rom[  946] = 'h00000050; 	    d_addr_rom[  946] = 'h00000f50; 	    wdata_rom[  946] = 'h922f6ba0; 	    wvalid_rom[  946] = 1; 
    i_addr_rom[  947] = 'h000007f0; 	    d_addr_rom[  947] = 'h00000c94; 	    wdata_rom[  947] = 'hcb193b58; 	    wvalid_rom[  947] = 0; 
    i_addr_rom[  948] = 'h00000784; 	    d_addr_rom[  948] = 'h00000e10; 	    wdata_rom[  948] = 'h0e99829e; 	    wvalid_rom[  948] = 1; 
    i_addr_rom[  949] = 'h000007c4; 	    d_addr_rom[  949] = 'h00000e34; 	    wdata_rom[  949] = 'h8349c51d; 	    wvalid_rom[  949] = 0; 
    i_addr_rom[  950] = 'h00000154; 	    d_addr_rom[  950] = 'h00000bf0; 	    wdata_rom[  950] = 'hdbcc7bca; 	    wvalid_rom[  950] = 0; 
    i_addr_rom[  951] = 'h00000408; 	    d_addr_rom[  951] = 'h00000a54; 	    wdata_rom[  951] = 'h6f1bae2f; 	    wvalid_rom[  951] = 0; 
    i_addr_rom[  952] = 'h0000066c; 	    d_addr_rom[  952] = 'h00000e20; 	    wdata_rom[  952] = 'hb610eac3; 	    wvalid_rom[  952] = 0; 
    i_addr_rom[  953] = 'h00000178; 	    d_addr_rom[  953] = 'h00000cf0; 	    wdata_rom[  953] = 'hf8cd501b; 	    wvalid_rom[  953] = 0; 
    i_addr_rom[  954] = 'h00000048; 	    d_addr_rom[  954] = 'h000008f4; 	    wdata_rom[  954] = 'h8e9e96ae; 	    wvalid_rom[  954] = 0; 
    i_addr_rom[  955] = 'h00000648; 	    d_addr_rom[  955] = 'h00000e9c; 	    wdata_rom[  955] = 'hff1f81bf; 	    wvalid_rom[  955] = 1; 
    i_addr_rom[  956] = 'h000000cc; 	    d_addr_rom[  956] = 'h000009b8; 	    wdata_rom[  956] = 'h9320bdb9; 	    wvalid_rom[  956] = 0; 
    i_addr_rom[  957] = 'h00000564; 	    d_addr_rom[  957] = 'h000009d0; 	    wdata_rom[  957] = 'h0025755f; 	    wvalid_rom[  957] = 1; 
    i_addr_rom[  958] = 'h000004bc; 	    d_addr_rom[  958] = 'h00000c98; 	    wdata_rom[  958] = 'h6ebcf10c; 	    wvalid_rom[  958] = 1; 
    i_addr_rom[  959] = 'h00000088; 	    d_addr_rom[  959] = 'h00000fc8; 	    wdata_rom[  959] = 'h652bc8ba; 	    wvalid_rom[  959] = 1; 
    i_addr_rom[  960] = 'h0000064c; 	    d_addr_rom[  960] = 'h00000b78; 	    wdata_rom[  960] = 'h0c5279f6; 	    wvalid_rom[  960] = 1; 
    i_addr_rom[  961] = 'h00000240; 	    d_addr_rom[  961] = 'h00000f48; 	    wdata_rom[  961] = 'h69e015d5; 	    wvalid_rom[  961] = 1; 
    i_addr_rom[  962] = 'h00000280; 	    d_addr_rom[  962] = 'h00000cd4; 	    wdata_rom[  962] = 'h489fe383; 	    wvalid_rom[  962] = 0; 
    i_addr_rom[  963] = 'h000002c4; 	    d_addr_rom[  963] = 'h000008ec; 	    wdata_rom[  963] = 'h36f108e9; 	    wvalid_rom[  963] = 1; 
    i_addr_rom[  964] = 'h00000764; 	    d_addr_rom[  964] = 'h00000820; 	    wdata_rom[  964] = 'h9716c468; 	    wvalid_rom[  964] = 0; 
    i_addr_rom[  965] = 'h0000053c; 	    d_addr_rom[  965] = 'h00000dcc; 	    wdata_rom[  965] = 'h6d767290; 	    wvalid_rom[  965] = 0; 
    i_addr_rom[  966] = 'h0000035c; 	    d_addr_rom[  966] = 'h00000ea0; 	    wdata_rom[  966] = 'hbd530b97; 	    wvalid_rom[  966] = 1; 
    i_addr_rom[  967] = 'h000000d0; 	    d_addr_rom[  967] = 'h00000b68; 	    wdata_rom[  967] = 'h37e8b7b6; 	    wvalid_rom[  967] = 1; 
    i_addr_rom[  968] = 'h00000538; 	    d_addr_rom[  968] = 'h00000b94; 	    wdata_rom[  968] = 'hed6f1334; 	    wvalid_rom[  968] = 0; 
    i_addr_rom[  969] = 'h00000630; 	    d_addr_rom[  969] = 'h00000c6c; 	    wdata_rom[  969] = 'h1e7778dc; 	    wvalid_rom[  969] = 0; 
    i_addr_rom[  970] = 'h0000045c; 	    d_addr_rom[  970] = 'h00000980; 	    wdata_rom[  970] = 'h0899badf; 	    wvalid_rom[  970] = 1; 
    i_addr_rom[  971] = 'h0000010c; 	    d_addr_rom[  971] = 'h000008fc; 	    wdata_rom[  971] = 'hbe6aa6c5; 	    wvalid_rom[  971] = 0; 
    i_addr_rom[  972] = 'h00000268; 	    d_addr_rom[  972] = 'h0000087c; 	    wdata_rom[  972] = 'h0f75d091; 	    wvalid_rom[  972] = 0; 
    i_addr_rom[  973] = 'h00000218; 	    d_addr_rom[  973] = 'h00000c14; 	    wdata_rom[  973] = 'h216cd04e; 	    wvalid_rom[  973] = 1; 
    i_addr_rom[  974] = 'h00000430; 	    d_addr_rom[  974] = 'h00000ad4; 	    wdata_rom[  974] = 'h026487ca; 	    wvalid_rom[  974] = 1; 
    i_addr_rom[  975] = 'h00000660; 	    d_addr_rom[  975] = 'h00000a38; 	    wdata_rom[  975] = 'hdb71756b; 	    wvalid_rom[  975] = 0; 
    i_addr_rom[  976] = 'h000005c8; 	    d_addr_rom[  976] = 'h00000d7c; 	    wdata_rom[  976] = 'h3c4278f5; 	    wvalid_rom[  976] = 1; 
    i_addr_rom[  977] = 'h000007a8; 	    d_addr_rom[  977] = 'h0000080c; 	    wdata_rom[  977] = 'h1f941992; 	    wvalid_rom[  977] = 0; 
    i_addr_rom[  978] = 'h0000004c; 	    d_addr_rom[  978] = 'h00000b6c; 	    wdata_rom[  978] = 'hc4f7ba40; 	    wvalid_rom[  978] = 0; 
    i_addr_rom[  979] = 'h000000ec; 	    d_addr_rom[  979] = 'h000008b0; 	    wdata_rom[  979] = 'h56a98895; 	    wvalid_rom[  979] = 0; 
    i_addr_rom[  980] = 'h000001ac; 	    d_addr_rom[  980] = 'h00000ae4; 	    wdata_rom[  980] = 'h32116e77; 	    wvalid_rom[  980] = 1; 
    i_addr_rom[  981] = 'h00000718; 	    d_addr_rom[  981] = 'h00000834; 	    wdata_rom[  981] = 'h8a3575e5; 	    wvalid_rom[  981] = 1; 
    i_addr_rom[  982] = 'h000004dc; 	    d_addr_rom[  982] = 'h00000e8c; 	    wdata_rom[  982] = 'h7bbdc40f; 	    wvalid_rom[  982] = 1; 
    i_addr_rom[  983] = 'h000003a4; 	    d_addr_rom[  983] = 'h00000ca0; 	    wdata_rom[  983] = 'h9a4bc642; 	    wvalid_rom[  983] = 0; 
    i_addr_rom[  984] = 'h000005a4; 	    d_addr_rom[  984] = 'h00000ea8; 	    wdata_rom[  984] = 'h4cf5e9a6; 	    wvalid_rom[  984] = 0; 
    i_addr_rom[  985] = 'h00000228; 	    d_addr_rom[  985] = 'h00000e88; 	    wdata_rom[  985] = 'h4152567a; 	    wvalid_rom[  985] = 1; 
    i_addr_rom[  986] = 'h00000248; 	    d_addr_rom[  986] = 'h0000087c; 	    wdata_rom[  986] = 'he6839600; 	    wvalid_rom[  986] = 0; 
    i_addr_rom[  987] = 'h00000690; 	    d_addr_rom[  987] = 'h00000fcc; 	    wdata_rom[  987] = 'h5c546645; 	    wvalid_rom[  987] = 0; 
    i_addr_rom[  988] = 'h00000358; 	    d_addr_rom[  988] = 'h000008dc; 	    wdata_rom[  988] = 'hd53fd327; 	    wvalid_rom[  988] = 1; 
    i_addr_rom[  989] = 'h00000634; 	    d_addr_rom[  989] = 'h00000fd8; 	    wdata_rom[  989] = 'h094509d7; 	    wvalid_rom[  989] = 1; 
    i_addr_rom[  990] = 'h00000008; 	    d_addr_rom[  990] = 'h00000f1c; 	    wdata_rom[  990] = 'hb1d07914; 	    wvalid_rom[  990] = 1; 
    i_addr_rom[  991] = 'h00000064; 	    d_addr_rom[  991] = 'h00000870; 	    wdata_rom[  991] = 'h70413197; 	    wvalid_rom[  991] = 1; 
    i_addr_rom[  992] = 'h000000f8; 	    d_addr_rom[  992] = 'h00000e70; 	    wdata_rom[  992] = 'hd0a57502; 	    wvalid_rom[  992] = 0; 
    i_addr_rom[  993] = 'h00000334; 	    d_addr_rom[  993] = 'h00000bc0; 	    wdata_rom[  993] = 'h8257dd08; 	    wvalid_rom[  993] = 1; 
    i_addr_rom[  994] = 'h000000e0; 	    d_addr_rom[  994] = 'h000009e0; 	    wdata_rom[  994] = 'h69258431; 	    wvalid_rom[  994] = 1; 
    i_addr_rom[  995] = 'h00000570; 	    d_addr_rom[  995] = 'h00000e04; 	    wdata_rom[  995] = 'hfba74cee; 	    wvalid_rom[  995] = 1; 
    i_addr_rom[  996] = 'h00000290; 	    d_addr_rom[  996] = 'h00000aac; 	    wdata_rom[  996] = 'h1313eed9; 	    wvalid_rom[  996] = 1; 
    i_addr_rom[  997] = 'h000007d0; 	    d_addr_rom[  997] = 'h00000ccc; 	    wdata_rom[  997] = 'h2c7703bd; 	    wvalid_rom[  997] = 1; 
    i_addr_rom[  998] = 'h000006a4; 	    d_addr_rom[  998] = 'h00000d84; 	    wdata_rom[  998] = 'h035eb9ad; 	    wvalid_rom[  998] = 1; 
    i_addr_rom[  999] = 'h000003d0; 	    d_addr_rom[  999] = 'h00000c3c; 	    wdata_rom[  999] = 'h8333cfcb; 	    wvalid_rom[  999] = 1; 
    i_addr_rom[ 1000] = 'h00000700; 	    d_addr_rom[ 1000] = 'h00000cf8; 	    wdata_rom[ 1000] = 'h2412f8c5; 	    wvalid_rom[ 1000] = 1; 
    i_addr_rom[ 1001] = 'h00000290; 	    d_addr_rom[ 1001] = 'h00000ef8; 	    wdata_rom[ 1001] = 'hb499c4df; 	    wvalid_rom[ 1001] = 1; 
    i_addr_rom[ 1002] = 'h000000e4; 	    d_addr_rom[ 1002] = 'h00000f58; 	    wdata_rom[ 1002] = 'h123d9e37; 	    wvalid_rom[ 1002] = 0; 
    i_addr_rom[ 1003] = 'h00000598; 	    d_addr_rom[ 1003] = 'h00000c64; 	    wdata_rom[ 1003] = 'hc9497c44; 	    wvalid_rom[ 1003] = 1; 
    i_addr_rom[ 1004] = 'h0000078c; 	    d_addr_rom[ 1004] = 'h00000df4; 	    wdata_rom[ 1004] = 'h10e7f5db; 	    wvalid_rom[ 1004] = 1; 
    i_addr_rom[ 1005] = 'h000007ac; 	    d_addr_rom[ 1005] = 'h00000be8; 	    wdata_rom[ 1005] = 'h1b577687; 	    wvalid_rom[ 1005] = 0; 
    i_addr_rom[ 1006] = 'h00000378; 	    d_addr_rom[ 1006] = 'h00000b24; 	    wdata_rom[ 1006] = 'h375d1324; 	    wvalid_rom[ 1006] = 0; 
    i_addr_rom[ 1007] = 'h00000050; 	    d_addr_rom[ 1007] = 'h00000c20; 	    wdata_rom[ 1007] = 'hbd981e5e; 	    wvalid_rom[ 1007] = 1; 
    i_addr_rom[ 1008] = 'h00000414; 	    d_addr_rom[ 1008] = 'h00000ac4; 	    wdata_rom[ 1008] = 'h81d59441; 	    wvalid_rom[ 1008] = 1; 
    i_addr_rom[ 1009] = 'h00000778; 	    d_addr_rom[ 1009] = 'h00000d88; 	    wdata_rom[ 1009] = 'h294fe69a; 	    wvalid_rom[ 1009] = 0; 
    i_addr_rom[ 1010] = 'h0000064c; 	    d_addr_rom[ 1010] = 'h000009d8; 	    wdata_rom[ 1010] = 'hecd681c0; 	    wvalid_rom[ 1010] = 1; 
    i_addr_rom[ 1011] = 'h00000110; 	    d_addr_rom[ 1011] = 'h00000c28; 	    wdata_rom[ 1011] = 'hd13021ac; 	    wvalid_rom[ 1011] = 0; 
    i_addr_rom[ 1012] = 'h00000130; 	    d_addr_rom[ 1012] = 'h00000fa8; 	    wdata_rom[ 1012] = 'h8dd9558e; 	    wvalid_rom[ 1012] = 1; 
    i_addr_rom[ 1013] = 'h000000b8; 	    d_addr_rom[ 1013] = 'h00000a5c; 	    wdata_rom[ 1013] = 'h7dd75454; 	    wvalid_rom[ 1013] = 1; 
    i_addr_rom[ 1014] = 'h00000698; 	    d_addr_rom[ 1014] = 'h000008c0; 	    wdata_rom[ 1014] = 'hc3db4ff7; 	    wvalid_rom[ 1014] = 0; 
    i_addr_rom[ 1015] = 'h000005fc; 	    d_addr_rom[ 1015] = 'h00000c9c; 	    wdata_rom[ 1015] = 'h7e9a41a0; 	    wvalid_rom[ 1015] = 1; 
    i_addr_rom[ 1016] = 'h000002bc; 	    d_addr_rom[ 1016] = 'h00000980; 	    wdata_rom[ 1016] = 'h9a9c30ba; 	    wvalid_rom[ 1016] = 1; 
    i_addr_rom[ 1017] = 'h000006b4; 	    d_addr_rom[ 1017] = 'h00000d6c; 	    wdata_rom[ 1017] = 'he57edc3b; 	    wvalid_rom[ 1017] = 0; 
    i_addr_rom[ 1018] = 'h00000394; 	    d_addr_rom[ 1018] = 'h00000f60; 	    wdata_rom[ 1018] = 'hd0412ccd; 	    wvalid_rom[ 1018] = 0; 
    i_addr_rom[ 1019] = 'h00000598; 	    d_addr_rom[ 1019] = 'h00000850; 	    wdata_rom[ 1019] = 'h0369638b; 	    wvalid_rom[ 1019] = 1; 
    i_addr_rom[ 1020] = 'h00000168; 	    d_addr_rom[ 1020] = 'h000009c8; 	    wdata_rom[ 1020] = 'h308f47fe; 	    wvalid_rom[ 1020] = 1; 
    i_addr_rom[ 1021] = 'h00000734; 	    d_addr_rom[ 1021] = 'h00000a34; 	    wdata_rom[ 1021] = 'h157cb48f; 	    wvalid_rom[ 1021] = 1; 
    i_addr_rom[ 1022] = 'h00000078; 	    d_addr_rom[ 1022] = 'h000009cc; 	    wdata_rom[ 1022] = 'he7964bc8; 	    wvalid_rom[ 1022] = 0; 
    i_addr_rom[ 1023] = 'h0000074c; 	    d_addr_rom[ 1023] = 'h00000f1c; 	    wdata_rom[ 1023] = 'hd65aa3f6; 	    wvalid_rom[ 1023] = 1; 

end
// for icache 
wire            i_rvalid_pipe;
wire            i_rready_pipe;
wire    [31:0]  i_raddr_pipe;
wire    [31:0]  i_rdata_pipe;
wire            i_rvalid;
wire            i_rready;
// icache && arbiter 
wire    [31:0]  i_raddr;
wire    [31:0]  i_rdata;
wire            i_rlast;
wire    [2:0]   i_rsize;
wire    [7:0]   i_rlen;
// icache_debug
reg             i_rvalid_ff;
reg     [31:0]  i_raddr_ff;
reg             i_error_reg;
reg             i_pass_reg;
wire    [31:0]  i_correct_data;

// for dcache
wire    [31:0]  d_addr_pipe;
wire            d_rvalid_pipe;
wire            d_rready_pipe;
wire    [31:0]  d_rdata_pipe;
wire            d_wvalid_pipe;
wire            d_wready_pipe;
wire    [31:0]  d_wdata_pipe;
wire    [3:0]   d_wstrb_pipe;
// dcache && arbiter
wire            d_rvalid;
wire            d_rready;
wire    [31:0]  d_raddr;
wire    [31:0]  d_rdata;
wire            d_rlast;
wire    [2:0]   d_rsize;
wire    [7:0]   d_rlen;
wire            d_wvalid;
wire            d_wready;
wire    [31:0]  d_waddr;
wire    [31:0]  d_wdata;
wire    [3:0]   d_wstrb;
wire            d_wlast;
wire    [2:0]   d_wsize;
wire    [7:0]   d_wlen;
wire            d_bvalid;
wire            d_bready;
// dcache_debug
reg             d_rvalid_ff;
reg             d_wvalid_ff;
reg     [31:0]  d_wdata_ff;
reg     [31:0]  d_addr_ff;
reg             d_error_reg;
reg             d_pass_reg;
wire    [31:0]  d_correct_data;

// arbiter with main mem
wire    [31:0]  araddr;
wire            arvalid;
wire            arready;
wire    [7:0]   arlen;
wire    [2:0]   arsize;
wire    [1:0]   arburst;
wire    [31:0]  rdata;
wire    [1:0]   rresp;
wire            rvalid;
wire            rready;
wire            rlast;
wire    [31:0]  awaddr;
wire            awvalid;
wire            awready;
wire    [7:0]   awlen;
wire    [2:0]   awsize;
wire    [1:0]   awburst;
wire    [31:0]  wdata;
wire    [3:0]   wstrb;
wire            wvalid;
wire            wready;
wire            wlast;
wire    [1:0]   bresp;
wire            bvalid;
wire            bready;

assign i_raddr_pipe = i_addr_rom[i_test_index];
assign i_correct_data = data_ram[i_raddr_ff >> 2];
assign i_rvalid_pipe = 1'b1;
// simulate IF1-IF2 register i_rvalid_ff && i_raddr_ff
always @(posedge clk) begin
    if(!rstn) begin
        i_rvalid_ff <= 0;
        i_raddr_ff <= 0;
    end
    else if(!(i_rvalid_ff && !i_rready_pipe))begin
        i_rvalid_ff <= i_rvalid_pipe;
        i_raddr_ff <= i_raddr_pipe;
    end
end
// update i_test_index
always @(posedge clk) begin
    if(!rstn) begin
        i_test_index <= 0;
        i_pass_reg <= 0;
    end
    else if (i_test_index >= (TOTAL_WORD_NUM / 2-1)) begin
        i_test_index <= (TOTAL_WORD_NUM / 2-1);
        i_pass_reg <= 1;
    end
    else if(!(i_rvalid_ff && !i_rready_pipe) && !i_error_reg) begin
        i_test_index <= i_test_index + 1;
    end
end
// update i_error 
always @(posedge clk) begin
    if(!rstn) begin
        i_error_reg <= 0;
    end
    else if(i_error_reg) begin
        i_error_reg <= 1;
    end
    else if(i_rvalid_ff && i_rready_pipe) begin
        i_error_reg <= !(i_rdata_pipe  == i_correct_data);
    end
end

assign d_addr_pipe           = d_addr_rom[d_test_index];
assign d_correct_data   = data_ram[d_addr_ff >> 2];
assign d_rvalid_pipe         = !wvalid_rom[d_test_index];
assign d_wvalid_pipe         = wvalid_rom[d_test_index];
assign d_wdata_pipe          = wdata_rom[d_test_index];
assign d_wstrb_pipe          = d_wvalid_pipe ? 4'b1111 : 4'b0000;
// simulate EX-MEM register
always @(posedge clk) begin
    if(!rstn) begin
        d_rvalid_ff <= 0;
        d_addr_ff   <= 0;
        d_wvalid_ff <= 0;
        d_wdata_ff  <= 0;
    end
    else if(!(d_rvalid_ff && !d_rready_pipe) && !(d_wvalid_ff && !d_wready_pipe))begin
        d_rvalid_ff <= d_rvalid_pipe;
        d_addr_ff   <= d_addr_pipe;
        d_wvalid_ff <= d_wvalid_pipe;
        d_wdata_ff  <= d_wdata_pipe;
    end
end
// update d_test_index
always @(posedge clk) begin
    if(!rstn) begin
        d_test_index    <= TOTAL_WORD_NUM / 2;
        d_pass_reg      <= 0;
    end
    else if (d_test_index >= (TOTAL_WORD_NUM-1)) begin
        d_test_index    <= (TOTAL_WORD_NUM-1);
        d_pass_reg      <= 1;
    end
    else if(!(d_rvalid_ff && !d_rready_pipe)  && !(d_wvalid_ff && !d_wready_pipe) && !d_error_reg) begin
        d_test_index    <= d_test_index + 1;
    end
end
// update data_ram
always @(posedge clk) begin
    if(d_wvalid_ff && d_wready_pipe) begin
        data_ram[d_addr_ff >> 2] <= d_wdata_ff;
    end
end
// update d_error 
always @(posedge clk) begin
    if(!rstn) begin
        d_error_reg <= 0;
    end
    else if(d_error_reg) begin
        d_error_reg <= 1;
    end
    else if(d_rvalid_ff && d_rready_pipe) begin
        d_error_reg <= !(d_rdata_pipe  == d_correct_data);
    end
end

icache #(
  .INDEX_WIDTH          (INDEX_WIDTH),
  .WORD_OFFSET_WIDTH    (WORD_OFFSET_WIDTH)
)
icache_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .rvalid   (i_rvalid_pipe ),
    .rready   (i_rready_pipe ),
    .raddr    (i_raddr_pipe ),
    .rdata    (i_rdata_pipe ),

    .i_rvalid (i_rvalid ),
    .i_rready (i_rready ),
    .i_raddr  (i_raddr ),
    .i_rdata  (i_rdata ),
    .i_rlast  (i_rlast ),
    .i_rsize  (i_rsize ),
    .i_rlen   (i_rlen)
);
dcache #(
    .INDEX_WIDTH        (INDEX_WIDTH ),
    .WORD_OFFSET_WIDTH  (WORD_OFFSET_WIDTH )
)
dcache_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .addr     (d_addr_pipe ),
    .rvalid   (d_rvalid_pipe ),
    .rready   (d_rready_pipe ),
    .rdata    (d_rdata_pipe ),
    .wvalid   (d_wvalid_pipe ),
    .wready   (d_wready_pipe ),
    .wdata    (d_wdata_pipe ),
    .wstrb    (d_wstrb_pipe ),
    .d_rvalid (d_rvalid ),
    .d_rready (d_rready ),
    .d_raddr  (d_raddr ),
    .d_rdata  (d_rdata ),
    .d_rlast  (d_rlast ),
    .d_rsize  (d_rsize ),
    .d_rlen   (d_rlen ),
    .d_wvalid (d_wvalid ),
    .d_wready (d_wready ),
    .d_waddr  (d_waddr ),
    .d_wdata  (d_wdata ),
    .d_wstrb  (d_wstrb ),
    .d_wlast  (d_wlast ),
    .d_wsize  (d_wsize ),
    .d_wlen   (d_wlen ),
    .d_bvalid (d_bvalid ),
    .d_bready (d_bready )
);

axi_arbiter axi_arbiter_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .i_rvalid (i_rvalid ),
    .i_rready (i_rready ),
    .i_raddr  (i_raddr ),
    .i_rdata  (i_rdata ),
    .i_rlast  (i_rlast ),
    .i_rsize  (i_rsize ),
    .i_rlen   (i_rlen ),
    .d_rvalid (d_rvalid ),
    .d_rready (d_rready ),
    .d_raddr  (d_raddr ),
    .d_rdata  (d_rdata ),
    .d_rlast  (d_rlast ),
    .d_rsize  (d_rsize ),
    .d_rlen   (d_rlen ),
    .d_wvalid (d_wvalid ),
    .d_wready (d_wready ),
    .d_waddr  (d_waddr ),
    .d_wdata  (d_wdata ),
    .d_wstrb  (d_wstrb ),
    .d_wlast  (d_wlast ),
    .d_wsize  (d_wsize ),
    .d_wlen   (d_wlen ),
    .d_bvalid (d_bvalid ),
    .d_bready (d_bready ),
    .araddr   (araddr ),
    .arvalid  (arvalid ),
    .arready  (arready ),
    .arlen    (arlen ),
    .arsize   (arsize ),
    .arburst  (arburst ),
    .rdata    (rdata ),
    .rresp    (rresp ),
    .rvalid   (rvalid ),
    .rready   (rready ),
    .rlast    (rlast ),
    .awaddr   (awaddr ),
    .awvalid  (awvalid ),
    .awready  (awready ),
    .awlen    (awlen ),
    .awsize   (awsize ),
    .awburst  (awburst ),
    .wdata    (wdata ),
    .wstrb    (wstrb ),
    .wvalid   (wvalid ),
    .wready   (wready ),
    .wlast    (wlast ),
    .bresp    (bresp ),
    .bvalid   (bvalid ),
    .bready   (bready)
);
main_memory main_mem(
    .s_aclk         (clk ),
    .s_aresetn      (rstn ),
    .s_axi_araddr   (araddr ),
    .s_axi_arburst  (arburst ),
    .s_axi_arid     (4'b0),
    .s_axi_arlen    (arlen ),
    .s_axi_arready  (arready ),
    .s_axi_arsize   (arsize ),
    .s_axi_arvalid  (arvalid ),
    .s_axi_awaddr   (awaddr ),
    .s_axi_awburst  (awburst ),
    .s_axi_awid     (4'b0),
    .s_axi_awlen    (awlen ),
    .s_axi_awready  (awready ),
    .s_axi_awsize   (awsize ),
    .s_axi_awvalid  (awvalid ),
    .s_axi_bid      (),
    .s_axi_bready   (bready ),
    .s_axi_bresp    (bresp ),
    .s_axi_bvalid   (bvalid ),
    .s_axi_rdata    (rdata ),
    .s_axi_rid      (),
    .s_axi_rlast    (rlast ),
    .s_axi_rready   (rready ),
    .s_axi_rresp    (rresp ),
    .s_axi_rvalid   (rvalid ),
    .s_axi_wdata    (wdata ),
    .s_axi_wlast    (wlast ),
    .s_axi_wready   (wready ),
    .s_axi_wstrb    (wstrb ),
    .s_axi_wvalid   (wvalid )
);
endmodule

